VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DSP48
  CLASS BLOCK ;
  FOREIGN DSP48 ;
  ORIGIN 0.000 0.000 ;
  SIZE 597.400 BY 600.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.400 596.000 1.680 600.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.800 596.000 158.080 600.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.440 596.000 173.720 600.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.080 596.000 189.360 600.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.720 596.000 205.000 600.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.360 596.000 220.640 600.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.000 596.000 236.280 600.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.640 596.000 251.920 600.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.280 596.000 267.560 600.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.920 596.000 283.200 600.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.560 596.000 298.840 600.000 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.040 596.000 17.320 600.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.200 596.000 314.480 600.000 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.840 596.000 330.120 600.000 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.480 596.000 345.760 600.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.120 596.000 361.400 600.000 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.760 596.000 377.040 600.000 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.400 596.000 392.680 600.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.040 596.000 408.320 600.000 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.680 596.000 423.960 600.000 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.320 596.000 439.600 600.000 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.960 596.000 455.240 600.000 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.680 596.000 32.960 600.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.600 596.000 470.880 600.000 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.240 596.000 486.520 600.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.880 596.000 502.160 600.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.520 596.000 517.800 600.000 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.160 596.000 533.440 600.000 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.800 596.000 549.080 600.000 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.440 596.000 564.720 600.000 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.080 596.000 580.360 600.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.320 596.000 48.600 600.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.960 596.000 64.240 600.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.600 596.000 79.880 600.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.240 596.000 95.520 600.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.880 596.000 111.160 600.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.520 596.000 126.800 600.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.160 596.000 142.440 600.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.460 596.000 6.740 600.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.860 596.000 163.140 600.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.500 596.000 178.780 600.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.140 596.000 194.420 600.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.780 596.000 210.060 600.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.420 596.000 225.700 600.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.060 596.000 241.340 600.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.700 596.000 256.980 600.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.340 596.000 272.620 600.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.980 596.000 288.260 600.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.620 596.000 303.900 600.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.100 596.000 22.380 600.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.260 596.000 319.540 600.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.900 596.000 335.180 600.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.540 596.000 350.820 600.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.180 596.000 366.460 600.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.820 596.000 382.100 600.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.460 596.000 397.740 600.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.100 596.000 413.380 600.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.740 596.000 429.020 600.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.380 596.000 444.660 600.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.020 596.000 460.300 600.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.740 596.000 38.020 600.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.660 596.000 475.940 600.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.300 596.000 491.580 600.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.940 596.000 507.220 600.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.580 596.000 522.860 600.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.220 596.000 538.500 600.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.860 596.000 554.140 600.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.500 596.000 569.780 600.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.140 596.000 585.420 600.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.380 596.000 53.660 600.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.020 596.000 69.300 600.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.660 596.000 84.940 600.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.300 596.000 100.580 600.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.940 596.000 116.220 600.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.580 596.000 131.860 600.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.220 596.000 147.500 600.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.520 596.000 11.800 600.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.920 596.000 168.200 600.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.560 596.000 183.840 600.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.200 596.000 199.480 600.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.840 596.000 215.120 600.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.480 596.000 230.760 600.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.120 596.000 246.400 600.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.760 596.000 262.040 600.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.400 596.000 277.680 600.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.040 596.000 293.320 600.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.140 596.000 309.420 600.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.160 596.000 27.440 600.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.780 596.000 325.060 600.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.420 596.000 340.700 600.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.060 596.000 356.340 600.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.700 596.000 371.980 600.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 387.340 596.000 387.620 600.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.980 596.000 403.260 600.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.620 596.000 418.900 600.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.260 596.000 434.540 600.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.900 596.000 450.180 600.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.540 596.000 465.820 600.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.800 596.000 43.080 600.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.180 596.000 481.460 600.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.820 596.000 497.100 600.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.460 596.000 512.740 600.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.100 596.000 528.380 600.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.740 596.000 544.020 600.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.380 596.000 559.660 600.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.020 596.000 575.300 600.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.660 596.000 590.940 600.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.440 596.000 58.720 600.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.080 596.000 74.360 600.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.720 596.000 90.000 600.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.360 596.000 105.640 600.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.000 596.000 121.280 600.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.640 596.000 136.920 600.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.280 596.000 152.560 600.000 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.280 0.000 267.560 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.720 0.000 527.000 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.480 0.000 529.760 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.240 0.000 532.520 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.540 0.000 534.820 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.300 0.000 537.580 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.060 0.000 540.340 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.360 0.000 542.640 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.120 0.000 545.400 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.880 0.000 548.160 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.180 0.000 550.460 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.040 0.000 293.320 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.940 0.000 553.220 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.700 0.000 555.980 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.000 0.000 558.280 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.760 0.000 561.040 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.060 0.000 563.340 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.820 0.000 566.100 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.580 0.000 568.860 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.880 0.000 571.160 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.640 0.000 573.920 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.400 0.000 576.680 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.800 0.000 296.080 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.700 0.000 578.980 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.460 0.000 581.740 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.220 0.000 584.500 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.520 0.000 586.800 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.280 0.000 589.560 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.040 0.000 592.320 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.340 0.000 594.620 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.100 0.000 597.380 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.560 0.000 298.840 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.860 0.000 301.140 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.620 0.000 303.900 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.380 0.000 306.660 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.680 0.000 308.960 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.440 0.000 311.720 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.200 0.000 314.480 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.500 0.000 316.780 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.040 0.000 270.320 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.260 0.000 319.540 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.560 0.000 321.840 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.320 0.000 324.600 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.080 0.000 327.360 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.380 0.000 329.660 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.140 0.000 332.420 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.900 0.000 335.180 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.200 0.000 337.480 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.960 0.000 340.240 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.720 0.000 343.000 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.340 0.000 272.620 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.020 0.000 345.300 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.780 0.000 348.060 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.540 0.000 350.820 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.840 0.000 353.120 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.600 0.000 355.880 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.360 0.000 358.640 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.660 0.000 360.940 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.420 0.000 363.700 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.720 0.000 366.000 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.480 0.000 368.760 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.100 0.000 275.380 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.240 0.000 371.520 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.540 0.000 373.820 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.300 0.000 376.580 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.060 0.000 379.340 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.360 0.000 381.640 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 384.120 0.000 384.400 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.880 0.000 387.160 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.180 0.000 389.460 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.940 0.000 392.220 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.700 0.000 394.980 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.860 0.000 278.140 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.000 0.000 397.280 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.760 0.000 400.040 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.060 0.000 402.340 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.820 0.000 405.100 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.580 0.000 407.860 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.880 0.000 410.160 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.640 0.000 412.920 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.400 0.000 415.680 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.700 0.000 417.980 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.460 0.000 420.740 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.160 0.000 280.440 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.220 0.000 423.500 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.520 0.000 425.800 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.280 0.000 428.560 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.040 0.000 431.320 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.340 0.000 433.620 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.100 0.000 436.380 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.860 0.000 439.140 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.160 0.000 441.440 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.920 0.000 444.200 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.220 0.000 446.500 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.920 0.000 283.200 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.980 0.000 449.260 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.740 0.000 452.020 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.040 0.000 454.320 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.800 0.000 457.080 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.560 0.000 459.840 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.860 0.000 462.140 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 464.620 0.000 464.900 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.380 0.000 467.660 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.680 0.000 469.960 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.440 0.000 472.720 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.220 0.000 285.500 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.200 0.000 475.480 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.500 0.000 477.780 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.260 0.000 480.540 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.560 0.000 482.840 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.320 0.000 485.600 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.080 0.000 488.360 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.380 0.000 490.660 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.140 0.000 493.420 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.900 0.000 496.180 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.200 0.000 498.480 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.980 0.000 288.260 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 500.960 0.000 501.240 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.720 0.000 504.000 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.020 0.000 506.300 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.780 0.000 509.060 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.540 0.000 511.820 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.840 0.000 514.120 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.600 0.000 516.880 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 519.360 0.000 519.640 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.660 0.000 521.940 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.420 0.000 524.700 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.740 0.000 291.020 4.000 ;
    END
  END la_data_in[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.720 596.000 596.000 600.000 ;
    END
  END user_clock2
  PIN wb_ACK
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.020 0.000 0.300 4.000 ;
    END
  END wb_ACK
  PIN wb_ADR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.960 0.000 18.240 4.000 ;
    END
  END wb_ADR[0]
  PIN wb_ADR[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.700 0.000 95.980 4.000 ;
    END
  END wb_ADR[10]
  PIN wb_ADR[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.520 0.000 103.800 4.000 ;
    END
  END wb_ADR[11]
  PIN wb_ADR[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.340 0.000 111.620 4.000 ;
    END
  END wb_ADR[12]
  PIN wb_ADR[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.160 0.000 119.440 4.000 ;
    END
  END wb_ADR[13]
  PIN wb_ADR[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.980 0.000 127.260 4.000 ;
    END
  END wb_ADR[14]
  PIN wb_ADR[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.800 0.000 135.080 4.000 ;
    END
  END wb_ADR[15]
  PIN wb_ADR[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.620 0.000 142.900 4.000 ;
    END
  END wb_ADR[16]
  PIN wb_ADR[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.440 0.000 150.720 4.000 ;
    END
  END wb_ADR[17]
  PIN wb_ADR[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.260 0.000 158.540 4.000 ;
    END
  END wb_ADR[18]
  PIN wb_ADR[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.080 0.000 166.360 4.000 ;
    END
  END wb_ADR[19]
  PIN wb_ADR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.780 0.000 26.060 4.000 ;
    END
  END wb_ADR[1]
  PIN wb_ADR[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.900 0.000 174.180 4.000 ;
    END
  END wb_ADR[20]
  PIN wb_ADR[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.720 0.000 182.000 4.000 ;
    END
  END wb_ADR[21]
  PIN wb_ADR[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.540 0.000 189.820 4.000 ;
    END
  END wb_ADR[22]
  PIN wb_ADR[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.360 0.000 197.640 4.000 ;
    END
  END wb_ADR[23]
  PIN wb_ADR[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.720 0.000 205.000 4.000 ;
    END
  END wb_ADR[24]
  PIN wb_ADR[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.540 0.000 212.820 4.000 ;
    END
  END wb_ADR[25]
  PIN wb_ADR[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.360 0.000 220.640 4.000 ;
    END
  END wb_ADR[26]
  PIN wb_ADR[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.180 0.000 228.460 4.000 ;
    END
  END wb_ADR[27]
  PIN wb_ADR[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.000 0.000 236.280 4.000 ;
    END
  END wb_ADR[28]
  PIN wb_ADR[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.820 0.000 244.100 4.000 ;
    END
  END wb_ADR[29]
  PIN wb_ADR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.600 0.000 33.880 4.000 ;
    END
  END wb_ADR[2]
  PIN wb_ADR[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.640 0.000 251.920 4.000 ;
    END
  END wb_ADR[30]
  PIN wb_ADR[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.460 0.000 259.740 4.000 ;
    END
  END wb_ADR[31]
  PIN wb_ADR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.420 0.000 41.700 4.000 ;
    END
  END wb_ADR[3]
  PIN wb_ADR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.240 0.000 49.520 4.000 ;
    END
  END wb_ADR[4]
  PIN wb_ADR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 57.060 0.000 57.340 4.000 ;
    END
  END wb_ADR[5]
  PIN wb_ADR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.880 0.000 65.160 4.000 ;
    END
  END wb_ADR[6]
  PIN wb_ADR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.700 0.000 72.980 4.000 ;
    END
  END wb_ADR[7]
  PIN wb_ADR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.060 0.000 80.340 4.000 ;
    END
  END wb_ADR[8]
  PIN wb_ADR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.880 0.000 88.160 4.000 ;
    END
  END wb_ADR[9]
  PIN wb_CYC
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.320 0.000 2.600 4.000 ;
    END
  END wb_CYC
  PIN wb_DAT_MISO[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.720 0.000 21.000 4.000 ;
    END
  END wb_DAT_MISO[0]
  PIN wb_DAT_MISO[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.460 0.000 98.740 4.000 ;
    END
  END wb_DAT_MISO[10]
  PIN wb_DAT_MISO[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.280 0.000 106.560 4.000 ;
    END
  END wb_DAT_MISO[11]
  PIN wb_DAT_MISO[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.100 0.000 114.380 4.000 ;
    END
  END wb_DAT_MISO[12]
  PIN wb_DAT_MISO[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.920 0.000 122.200 4.000 ;
    END
  END wb_DAT_MISO[13]
  PIN wb_DAT_MISO[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.740 0.000 130.020 4.000 ;
    END
  END wb_DAT_MISO[14]
  PIN wb_DAT_MISO[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.560 0.000 137.840 4.000 ;
    END
  END wb_DAT_MISO[15]
  PIN wb_DAT_MISO[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.380 0.000 145.660 4.000 ;
    END
  END wb_DAT_MISO[16]
  PIN wb_DAT_MISO[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.200 0.000 153.480 4.000 ;
    END
  END wb_DAT_MISO[17]
  PIN wb_DAT_MISO[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.560 0.000 160.840 4.000 ;
    END
  END wb_DAT_MISO[18]
  PIN wb_DAT_MISO[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.380 0.000 168.660 4.000 ;
    END
  END wb_DAT_MISO[19]
  PIN wb_DAT_MISO[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.540 0.000 28.820 4.000 ;
    END
  END wb_DAT_MISO[1]
  PIN wb_DAT_MISO[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.200 0.000 176.480 4.000 ;
    END
  END wb_DAT_MISO[20]
  PIN wb_DAT_MISO[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.020 0.000 184.300 4.000 ;
    END
  END wb_DAT_MISO[21]
  PIN wb_DAT_MISO[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.840 0.000 192.120 4.000 ;
    END
  END wb_DAT_MISO[22]
  PIN wb_DAT_MISO[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.660 0.000 199.940 4.000 ;
    END
  END wb_DAT_MISO[23]
  PIN wb_DAT_MISO[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.480 0.000 207.760 4.000 ;
    END
  END wb_DAT_MISO[24]
  PIN wb_DAT_MISO[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.300 0.000 215.580 4.000 ;
    END
  END wb_DAT_MISO[25]
  PIN wb_DAT_MISO[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.120 0.000 223.400 4.000 ;
    END
  END wb_DAT_MISO[26]
  PIN wb_DAT_MISO[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.940 0.000 231.220 4.000 ;
    END
  END wb_DAT_MISO[27]
  PIN wb_DAT_MISO[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.760 0.000 239.040 4.000 ;
    END
  END wb_DAT_MISO[28]
  PIN wb_DAT_MISO[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.580 0.000 246.860 4.000 ;
    END
  END wb_DAT_MISO[29]
  PIN wb_DAT_MISO[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.360 0.000 36.640 4.000 ;
    END
  END wb_DAT_MISO[2]
  PIN wb_DAT_MISO[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.400 0.000 254.680 4.000 ;
    END
  END wb_DAT_MISO[30]
  PIN wb_DAT_MISO[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.220 0.000 262.500 4.000 ;
    END
  END wb_DAT_MISO[31]
  PIN wb_DAT_MISO[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.720 0.000 44.000 4.000 ;
    END
  END wb_DAT_MISO[3]
  PIN wb_DAT_MISO[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.540 0.000 51.820 4.000 ;
    END
  END wb_DAT_MISO[4]
  PIN wb_DAT_MISO[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.360 0.000 59.640 4.000 ;
    END
  END wb_DAT_MISO[5]
  PIN wb_DAT_MISO[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.180 0.000 67.460 4.000 ;
    END
  END wb_DAT_MISO[6]
  PIN wb_DAT_MISO[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.000 0.000 75.280 4.000 ;
    END
  END wb_DAT_MISO[7]
  PIN wb_DAT_MISO[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.820 0.000 83.100 4.000 ;
    END
  END wb_DAT_MISO[8]
  PIN wb_DAT_MISO[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.640 0.000 90.920 4.000 ;
    END
  END wb_DAT_MISO[9]
  PIN wb_DAT_MOSI[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.020 0.000 23.300 4.000 ;
    END
  END wb_DAT_MOSI[0]
  PIN wb_DAT_MOSI[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.220 0.000 101.500 4.000 ;
    END
  END wb_DAT_MOSI[10]
  PIN wb_DAT_MOSI[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.040 0.000 109.320 4.000 ;
    END
  END wb_DAT_MOSI[11]
  PIN wb_DAT_MOSI[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.860 0.000 117.140 4.000 ;
    END
  END wb_DAT_MOSI[12]
  PIN wb_DAT_MOSI[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.220 0.000 124.500 4.000 ;
    END
  END wb_DAT_MOSI[13]
  PIN wb_DAT_MOSI[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.040 0.000 132.320 4.000 ;
    END
  END wb_DAT_MOSI[14]
  PIN wb_DAT_MOSI[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.860 0.000 140.140 4.000 ;
    END
  END wb_DAT_MOSI[15]
  PIN wb_DAT_MOSI[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.680 0.000 147.960 4.000 ;
    END
  END wb_DAT_MOSI[16]
  PIN wb_DAT_MOSI[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.500 0.000 155.780 4.000 ;
    END
  END wb_DAT_MOSI[17]
  PIN wb_DAT_MOSI[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.320 0.000 163.600 4.000 ;
    END
  END wb_DAT_MOSI[18]
  PIN wb_DAT_MOSI[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.140 0.000 171.420 4.000 ;
    END
  END wb_DAT_MOSI[19]
  PIN wb_DAT_MOSI[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.840 0.000 31.120 4.000 ;
    END
  END wb_DAT_MOSI[1]
  PIN wb_DAT_MOSI[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.960 0.000 179.240 4.000 ;
    END
  END wb_DAT_MOSI[20]
  PIN wb_DAT_MOSI[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.780 0.000 187.060 4.000 ;
    END
  END wb_DAT_MOSI[21]
  PIN wb_DAT_MOSI[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.600 0.000 194.880 4.000 ;
    END
  END wb_DAT_MOSI[22]
  PIN wb_DAT_MOSI[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.420 0.000 202.700 4.000 ;
    END
  END wb_DAT_MOSI[23]
  PIN wb_DAT_MOSI[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.240 0.000 210.520 4.000 ;
    END
  END wb_DAT_MOSI[24]
  PIN wb_DAT_MOSI[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.060 0.000 218.340 4.000 ;
    END
  END wb_DAT_MOSI[25]
  PIN wb_DAT_MOSI[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.880 0.000 226.160 4.000 ;
    END
  END wb_DAT_MOSI[26]
  PIN wb_DAT_MOSI[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.700 0.000 233.980 4.000 ;
    END
  END wb_DAT_MOSI[27]
  PIN wb_DAT_MOSI[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.060 0.000 241.340 4.000 ;
    END
  END wb_DAT_MOSI[28]
  PIN wb_DAT_MOSI[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.880 0.000 249.160 4.000 ;
    END
  END wb_DAT_MOSI[29]
  PIN wb_DAT_MOSI[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.660 0.000 38.940 4.000 ;
    END
  END wb_DAT_MOSI[2]
  PIN wb_DAT_MOSI[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.700 0.000 256.980 4.000 ;
    END
  END wb_DAT_MOSI[30]
  PIN wb_DAT_MOSI[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.520 0.000 264.800 4.000 ;
    END
  END wb_DAT_MOSI[31]
  PIN wb_DAT_MOSI[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.480 0.000 46.760 4.000 ;
    END
  END wb_DAT_MOSI[3]
  PIN wb_DAT_MOSI[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.300 0.000 54.580 4.000 ;
    END
  END wb_DAT_MOSI[4]
  PIN wb_DAT_MOSI[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.120 0.000 62.400 4.000 ;
    END
  END wb_DAT_MOSI[5]
  PIN wb_DAT_MOSI[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.940 0.000 70.220 4.000 ;
    END
  END wb_DAT_MOSI[6]
  PIN wb_DAT_MOSI[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.760 0.000 78.040 4.000 ;
    END
  END wb_DAT_MOSI[7]
  PIN wb_DAT_MOSI[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.580 0.000 85.860 4.000 ;
    END
  END wb_DAT_MOSI[8]
  PIN wb_DAT_MOSI[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.400 0.000 93.680 4.000 ;
    END
  END wb_DAT_MOSI[9]
  PIN wb_SEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.080 0.000 5.360 4.000 ;
    END
  END wb_SEL
  PIN wb_STB
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.380 0.000 7.660 4.000 ;
    END
  END wb_STB
  PIN wb_WE
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.140 0.000 10.420 4.000 ;
    END
  END wb_WE
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.900 0.000 13.180 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.200 0.000 15.480 4.000 ;
    END
  END wb_rst_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 480.850 10.640 482.450 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 327.250 10.640 328.850 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 173.650 10.640 175.250 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 20.050 10.640 21.650 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 557.650 10.640 559.250 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 404.050 10.640 405.650 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 250.450 10.640 252.050 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 96.850 10.640 98.450 587.760 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 484.150 10.880 485.750 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 330.550 10.880 332.150 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 176.950 10.880 178.550 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 23.350 10.880 24.950 587.520 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 560.950 10.880 562.550 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 407.350 10.880 408.950 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 253.750 10.880 255.350 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 100.150 10.880 101.750 587.520 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 487.450 10.880 489.050 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 333.850 10.880 335.450 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 180.250 10.880 181.850 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 26.650 10.880 28.250 587.520 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 564.250 10.880 565.850 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 410.650 10.880 412.250 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 257.050 10.880 258.650 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 103.450 10.880 105.050 587.520 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 490.750 10.880 492.350 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 337.150 10.880 338.750 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 183.550 10.880 185.150 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 29.950 10.880 31.550 587.520 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 567.550 10.880 569.150 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 413.950 10.880 415.550 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 260.350 10.880 261.950 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 106.750 10.880 108.350 587.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 4.530 10.795 593.330 587.605 ;
      LAYER met1 ;
        RECT 0.000 4.460 597.400 587.760 ;
      LAYER met2 ;
        RECT 0.030 595.720 1.120 596.000 ;
        RECT 1.960 595.720 6.180 596.000 ;
        RECT 7.020 595.720 11.240 596.000 ;
        RECT 12.080 595.720 16.760 596.000 ;
        RECT 17.600 595.720 21.820 596.000 ;
        RECT 22.660 595.720 26.880 596.000 ;
        RECT 27.720 595.720 32.400 596.000 ;
        RECT 33.240 595.720 37.460 596.000 ;
        RECT 38.300 595.720 42.520 596.000 ;
        RECT 43.360 595.720 48.040 596.000 ;
        RECT 48.880 595.720 53.100 596.000 ;
        RECT 53.940 595.720 58.160 596.000 ;
        RECT 59.000 595.720 63.680 596.000 ;
        RECT 64.520 595.720 68.740 596.000 ;
        RECT 69.580 595.720 73.800 596.000 ;
        RECT 74.640 595.720 79.320 596.000 ;
        RECT 80.160 595.720 84.380 596.000 ;
        RECT 85.220 595.720 89.440 596.000 ;
        RECT 90.280 595.720 94.960 596.000 ;
        RECT 95.800 595.720 100.020 596.000 ;
        RECT 100.860 595.720 105.080 596.000 ;
        RECT 105.920 595.720 110.600 596.000 ;
        RECT 111.440 595.720 115.660 596.000 ;
        RECT 116.500 595.720 120.720 596.000 ;
        RECT 121.560 595.720 126.240 596.000 ;
        RECT 127.080 595.720 131.300 596.000 ;
        RECT 132.140 595.720 136.360 596.000 ;
        RECT 137.200 595.720 141.880 596.000 ;
        RECT 142.720 595.720 146.940 596.000 ;
        RECT 147.780 595.720 152.000 596.000 ;
        RECT 152.840 595.720 157.520 596.000 ;
        RECT 158.360 595.720 162.580 596.000 ;
        RECT 163.420 595.720 167.640 596.000 ;
        RECT 168.480 595.720 173.160 596.000 ;
        RECT 174.000 595.720 178.220 596.000 ;
        RECT 179.060 595.720 183.280 596.000 ;
        RECT 184.120 595.720 188.800 596.000 ;
        RECT 189.640 595.720 193.860 596.000 ;
        RECT 194.700 595.720 198.920 596.000 ;
        RECT 199.760 595.720 204.440 596.000 ;
        RECT 205.280 595.720 209.500 596.000 ;
        RECT 210.340 595.720 214.560 596.000 ;
        RECT 215.400 595.720 220.080 596.000 ;
        RECT 220.920 595.720 225.140 596.000 ;
        RECT 225.980 595.720 230.200 596.000 ;
        RECT 231.040 595.720 235.720 596.000 ;
        RECT 236.560 595.720 240.780 596.000 ;
        RECT 241.620 595.720 245.840 596.000 ;
        RECT 246.680 595.720 251.360 596.000 ;
        RECT 252.200 595.720 256.420 596.000 ;
        RECT 257.260 595.720 261.480 596.000 ;
        RECT 262.320 595.720 267.000 596.000 ;
        RECT 267.840 595.720 272.060 596.000 ;
        RECT 272.900 595.720 277.120 596.000 ;
        RECT 277.960 595.720 282.640 596.000 ;
        RECT 283.480 595.720 287.700 596.000 ;
        RECT 288.540 595.720 292.760 596.000 ;
        RECT 293.600 595.720 298.280 596.000 ;
        RECT 299.120 595.720 303.340 596.000 ;
        RECT 304.180 595.720 308.860 596.000 ;
        RECT 309.700 595.720 313.920 596.000 ;
        RECT 314.760 595.720 318.980 596.000 ;
        RECT 319.820 595.720 324.500 596.000 ;
        RECT 325.340 595.720 329.560 596.000 ;
        RECT 330.400 595.720 334.620 596.000 ;
        RECT 335.460 595.720 340.140 596.000 ;
        RECT 340.980 595.720 345.200 596.000 ;
        RECT 346.040 595.720 350.260 596.000 ;
        RECT 351.100 595.720 355.780 596.000 ;
        RECT 356.620 595.720 360.840 596.000 ;
        RECT 361.680 595.720 365.900 596.000 ;
        RECT 366.740 595.720 371.420 596.000 ;
        RECT 372.260 595.720 376.480 596.000 ;
        RECT 377.320 595.720 381.540 596.000 ;
        RECT 382.380 595.720 387.060 596.000 ;
        RECT 387.900 595.720 392.120 596.000 ;
        RECT 392.960 595.720 397.180 596.000 ;
        RECT 398.020 595.720 402.700 596.000 ;
        RECT 403.540 595.720 407.760 596.000 ;
        RECT 408.600 595.720 412.820 596.000 ;
        RECT 413.660 595.720 418.340 596.000 ;
        RECT 419.180 595.720 423.400 596.000 ;
        RECT 424.240 595.720 428.460 596.000 ;
        RECT 429.300 595.720 433.980 596.000 ;
        RECT 434.820 595.720 439.040 596.000 ;
        RECT 439.880 595.720 444.100 596.000 ;
        RECT 444.940 595.720 449.620 596.000 ;
        RECT 450.460 595.720 454.680 596.000 ;
        RECT 455.520 595.720 459.740 596.000 ;
        RECT 460.580 595.720 465.260 596.000 ;
        RECT 466.100 595.720 470.320 596.000 ;
        RECT 471.160 595.720 475.380 596.000 ;
        RECT 476.220 595.720 480.900 596.000 ;
        RECT 481.740 595.720 485.960 596.000 ;
        RECT 486.800 595.720 491.020 596.000 ;
        RECT 491.860 595.720 496.540 596.000 ;
        RECT 497.380 595.720 501.600 596.000 ;
        RECT 502.440 595.720 506.660 596.000 ;
        RECT 507.500 595.720 512.180 596.000 ;
        RECT 513.020 595.720 517.240 596.000 ;
        RECT 518.080 595.720 522.300 596.000 ;
        RECT 523.140 595.720 527.820 596.000 ;
        RECT 528.660 595.720 532.880 596.000 ;
        RECT 533.720 595.720 537.940 596.000 ;
        RECT 538.780 595.720 543.460 596.000 ;
        RECT 544.300 595.720 548.520 596.000 ;
        RECT 549.360 595.720 553.580 596.000 ;
        RECT 554.420 595.720 559.100 596.000 ;
        RECT 559.940 595.720 564.160 596.000 ;
        RECT 565.000 595.720 569.220 596.000 ;
        RECT 570.060 595.720 574.740 596.000 ;
        RECT 575.580 595.720 579.800 596.000 ;
        RECT 580.640 595.720 584.860 596.000 ;
        RECT 585.700 595.720 590.380 596.000 ;
        RECT 591.220 595.720 595.440 596.000 ;
        RECT 596.280 595.720 597.370 596.000 ;
        RECT 0.030 4.280 597.370 595.720 ;
        RECT 0.580 4.000 2.040 4.280 ;
        RECT 2.880 4.000 4.800 4.280 ;
        RECT 5.640 4.000 7.100 4.280 ;
        RECT 7.940 4.000 9.860 4.280 ;
        RECT 10.700 4.000 12.620 4.280 ;
        RECT 13.460 4.000 14.920 4.280 ;
        RECT 15.760 4.000 17.680 4.280 ;
        RECT 18.520 4.000 20.440 4.280 ;
        RECT 21.280 4.000 22.740 4.280 ;
        RECT 23.580 4.000 25.500 4.280 ;
        RECT 26.340 4.000 28.260 4.280 ;
        RECT 29.100 4.000 30.560 4.280 ;
        RECT 31.400 4.000 33.320 4.280 ;
        RECT 34.160 4.000 36.080 4.280 ;
        RECT 36.920 4.000 38.380 4.280 ;
        RECT 39.220 4.000 41.140 4.280 ;
        RECT 41.980 4.000 43.440 4.280 ;
        RECT 44.280 4.000 46.200 4.280 ;
        RECT 47.040 4.000 48.960 4.280 ;
        RECT 49.800 4.000 51.260 4.280 ;
        RECT 52.100 4.000 54.020 4.280 ;
        RECT 54.860 4.000 56.780 4.280 ;
        RECT 57.620 4.000 59.080 4.280 ;
        RECT 59.920 4.000 61.840 4.280 ;
        RECT 62.680 4.000 64.600 4.280 ;
        RECT 65.440 4.000 66.900 4.280 ;
        RECT 67.740 4.000 69.660 4.280 ;
        RECT 70.500 4.000 72.420 4.280 ;
        RECT 73.260 4.000 74.720 4.280 ;
        RECT 75.560 4.000 77.480 4.280 ;
        RECT 78.320 4.000 79.780 4.280 ;
        RECT 80.620 4.000 82.540 4.280 ;
        RECT 83.380 4.000 85.300 4.280 ;
        RECT 86.140 4.000 87.600 4.280 ;
        RECT 88.440 4.000 90.360 4.280 ;
        RECT 91.200 4.000 93.120 4.280 ;
        RECT 93.960 4.000 95.420 4.280 ;
        RECT 96.260 4.000 98.180 4.280 ;
        RECT 99.020 4.000 100.940 4.280 ;
        RECT 101.780 4.000 103.240 4.280 ;
        RECT 104.080 4.000 106.000 4.280 ;
        RECT 106.840 4.000 108.760 4.280 ;
        RECT 109.600 4.000 111.060 4.280 ;
        RECT 111.900 4.000 113.820 4.280 ;
        RECT 114.660 4.000 116.580 4.280 ;
        RECT 117.420 4.000 118.880 4.280 ;
        RECT 119.720 4.000 121.640 4.280 ;
        RECT 122.480 4.000 123.940 4.280 ;
        RECT 124.780 4.000 126.700 4.280 ;
        RECT 127.540 4.000 129.460 4.280 ;
        RECT 130.300 4.000 131.760 4.280 ;
        RECT 132.600 4.000 134.520 4.280 ;
        RECT 135.360 4.000 137.280 4.280 ;
        RECT 138.120 4.000 139.580 4.280 ;
        RECT 140.420 4.000 142.340 4.280 ;
        RECT 143.180 4.000 145.100 4.280 ;
        RECT 145.940 4.000 147.400 4.280 ;
        RECT 148.240 4.000 150.160 4.280 ;
        RECT 151.000 4.000 152.920 4.280 ;
        RECT 153.760 4.000 155.220 4.280 ;
        RECT 156.060 4.000 157.980 4.280 ;
        RECT 158.820 4.000 160.280 4.280 ;
        RECT 161.120 4.000 163.040 4.280 ;
        RECT 163.880 4.000 165.800 4.280 ;
        RECT 166.640 4.000 168.100 4.280 ;
        RECT 168.940 4.000 170.860 4.280 ;
        RECT 171.700 4.000 173.620 4.280 ;
        RECT 174.460 4.000 175.920 4.280 ;
        RECT 176.760 4.000 178.680 4.280 ;
        RECT 179.520 4.000 181.440 4.280 ;
        RECT 182.280 4.000 183.740 4.280 ;
        RECT 184.580 4.000 186.500 4.280 ;
        RECT 187.340 4.000 189.260 4.280 ;
        RECT 190.100 4.000 191.560 4.280 ;
        RECT 192.400 4.000 194.320 4.280 ;
        RECT 195.160 4.000 197.080 4.280 ;
        RECT 197.920 4.000 199.380 4.280 ;
        RECT 200.220 4.000 202.140 4.280 ;
        RECT 202.980 4.000 204.440 4.280 ;
        RECT 205.280 4.000 207.200 4.280 ;
        RECT 208.040 4.000 209.960 4.280 ;
        RECT 210.800 4.000 212.260 4.280 ;
        RECT 213.100 4.000 215.020 4.280 ;
        RECT 215.860 4.000 217.780 4.280 ;
        RECT 218.620 4.000 220.080 4.280 ;
        RECT 220.920 4.000 222.840 4.280 ;
        RECT 223.680 4.000 225.600 4.280 ;
        RECT 226.440 4.000 227.900 4.280 ;
        RECT 228.740 4.000 230.660 4.280 ;
        RECT 231.500 4.000 233.420 4.280 ;
        RECT 234.260 4.000 235.720 4.280 ;
        RECT 236.560 4.000 238.480 4.280 ;
        RECT 239.320 4.000 240.780 4.280 ;
        RECT 241.620 4.000 243.540 4.280 ;
        RECT 244.380 4.000 246.300 4.280 ;
        RECT 247.140 4.000 248.600 4.280 ;
        RECT 249.440 4.000 251.360 4.280 ;
        RECT 252.200 4.000 254.120 4.280 ;
        RECT 254.960 4.000 256.420 4.280 ;
        RECT 257.260 4.000 259.180 4.280 ;
        RECT 260.020 4.000 261.940 4.280 ;
        RECT 262.780 4.000 264.240 4.280 ;
        RECT 265.080 4.000 267.000 4.280 ;
        RECT 267.840 4.000 269.760 4.280 ;
        RECT 270.600 4.000 272.060 4.280 ;
        RECT 272.900 4.000 274.820 4.280 ;
        RECT 275.660 4.000 277.580 4.280 ;
        RECT 278.420 4.000 279.880 4.280 ;
        RECT 280.720 4.000 282.640 4.280 ;
        RECT 283.480 4.000 284.940 4.280 ;
        RECT 285.780 4.000 287.700 4.280 ;
        RECT 288.540 4.000 290.460 4.280 ;
        RECT 291.300 4.000 292.760 4.280 ;
        RECT 293.600 4.000 295.520 4.280 ;
        RECT 296.360 4.000 298.280 4.280 ;
        RECT 299.120 4.000 300.580 4.280 ;
        RECT 301.420 4.000 303.340 4.280 ;
        RECT 304.180 4.000 306.100 4.280 ;
        RECT 306.940 4.000 308.400 4.280 ;
        RECT 309.240 4.000 311.160 4.280 ;
        RECT 312.000 4.000 313.920 4.280 ;
        RECT 314.760 4.000 316.220 4.280 ;
        RECT 317.060 4.000 318.980 4.280 ;
        RECT 319.820 4.000 321.280 4.280 ;
        RECT 322.120 4.000 324.040 4.280 ;
        RECT 324.880 4.000 326.800 4.280 ;
        RECT 327.640 4.000 329.100 4.280 ;
        RECT 329.940 4.000 331.860 4.280 ;
        RECT 332.700 4.000 334.620 4.280 ;
        RECT 335.460 4.000 336.920 4.280 ;
        RECT 337.760 4.000 339.680 4.280 ;
        RECT 340.520 4.000 342.440 4.280 ;
        RECT 343.280 4.000 344.740 4.280 ;
        RECT 345.580 4.000 347.500 4.280 ;
        RECT 348.340 4.000 350.260 4.280 ;
        RECT 351.100 4.000 352.560 4.280 ;
        RECT 353.400 4.000 355.320 4.280 ;
        RECT 356.160 4.000 358.080 4.280 ;
        RECT 358.920 4.000 360.380 4.280 ;
        RECT 361.220 4.000 363.140 4.280 ;
        RECT 363.980 4.000 365.440 4.280 ;
        RECT 366.280 4.000 368.200 4.280 ;
        RECT 369.040 4.000 370.960 4.280 ;
        RECT 371.800 4.000 373.260 4.280 ;
        RECT 374.100 4.000 376.020 4.280 ;
        RECT 376.860 4.000 378.780 4.280 ;
        RECT 379.620 4.000 381.080 4.280 ;
        RECT 381.920 4.000 383.840 4.280 ;
        RECT 384.680 4.000 386.600 4.280 ;
        RECT 387.440 4.000 388.900 4.280 ;
        RECT 389.740 4.000 391.660 4.280 ;
        RECT 392.500 4.000 394.420 4.280 ;
        RECT 395.260 4.000 396.720 4.280 ;
        RECT 397.560 4.000 399.480 4.280 ;
        RECT 400.320 4.000 401.780 4.280 ;
        RECT 402.620 4.000 404.540 4.280 ;
        RECT 405.380 4.000 407.300 4.280 ;
        RECT 408.140 4.000 409.600 4.280 ;
        RECT 410.440 4.000 412.360 4.280 ;
        RECT 413.200 4.000 415.120 4.280 ;
        RECT 415.960 4.000 417.420 4.280 ;
        RECT 418.260 4.000 420.180 4.280 ;
        RECT 421.020 4.000 422.940 4.280 ;
        RECT 423.780 4.000 425.240 4.280 ;
        RECT 426.080 4.000 428.000 4.280 ;
        RECT 428.840 4.000 430.760 4.280 ;
        RECT 431.600 4.000 433.060 4.280 ;
        RECT 433.900 4.000 435.820 4.280 ;
        RECT 436.660 4.000 438.580 4.280 ;
        RECT 439.420 4.000 440.880 4.280 ;
        RECT 441.720 4.000 443.640 4.280 ;
        RECT 444.480 4.000 445.940 4.280 ;
        RECT 446.780 4.000 448.700 4.280 ;
        RECT 449.540 4.000 451.460 4.280 ;
        RECT 452.300 4.000 453.760 4.280 ;
        RECT 454.600 4.000 456.520 4.280 ;
        RECT 457.360 4.000 459.280 4.280 ;
        RECT 460.120 4.000 461.580 4.280 ;
        RECT 462.420 4.000 464.340 4.280 ;
        RECT 465.180 4.000 467.100 4.280 ;
        RECT 467.940 4.000 469.400 4.280 ;
        RECT 470.240 4.000 472.160 4.280 ;
        RECT 473.000 4.000 474.920 4.280 ;
        RECT 475.760 4.000 477.220 4.280 ;
        RECT 478.060 4.000 479.980 4.280 ;
        RECT 480.820 4.000 482.280 4.280 ;
        RECT 483.120 4.000 485.040 4.280 ;
        RECT 485.880 4.000 487.800 4.280 ;
        RECT 488.640 4.000 490.100 4.280 ;
        RECT 490.940 4.000 492.860 4.280 ;
        RECT 493.700 4.000 495.620 4.280 ;
        RECT 496.460 4.000 497.920 4.280 ;
        RECT 498.760 4.000 500.680 4.280 ;
        RECT 501.520 4.000 503.440 4.280 ;
        RECT 504.280 4.000 505.740 4.280 ;
        RECT 506.580 4.000 508.500 4.280 ;
        RECT 509.340 4.000 511.260 4.280 ;
        RECT 512.100 4.000 513.560 4.280 ;
        RECT 514.400 4.000 516.320 4.280 ;
        RECT 517.160 4.000 519.080 4.280 ;
        RECT 519.920 4.000 521.380 4.280 ;
        RECT 522.220 4.000 524.140 4.280 ;
        RECT 524.980 4.000 526.440 4.280 ;
        RECT 527.280 4.000 529.200 4.280 ;
        RECT 530.040 4.000 531.960 4.280 ;
        RECT 532.800 4.000 534.260 4.280 ;
        RECT 535.100 4.000 537.020 4.280 ;
        RECT 537.860 4.000 539.780 4.280 ;
        RECT 540.620 4.000 542.080 4.280 ;
        RECT 542.920 4.000 544.840 4.280 ;
        RECT 545.680 4.000 547.600 4.280 ;
        RECT 548.440 4.000 549.900 4.280 ;
        RECT 550.740 4.000 552.660 4.280 ;
        RECT 553.500 4.000 555.420 4.280 ;
        RECT 556.260 4.000 557.720 4.280 ;
        RECT 558.560 4.000 560.480 4.280 ;
        RECT 561.320 4.000 562.780 4.280 ;
        RECT 563.620 4.000 565.540 4.280 ;
        RECT 566.380 4.000 568.300 4.280 ;
        RECT 569.140 4.000 570.600 4.280 ;
        RECT 571.440 4.000 573.360 4.280 ;
        RECT 574.200 4.000 576.120 4.280 ;
        RECT 576.960 4.000 578.420 4.280 ;
        RECT 579.260 4.000 581.180 4.280 ;
        RECT 582.020 4.000 583.940 4.280 ;
        RECT 584.780 4.000 586.240 4.280 ;
        RECT 587.080 4.000 589.000 4.280 ;
        RECT 589.840 4.000 591.760 4.280 ;
        RECT 592.600 4.000 594.060 4.280 ;
        RECT 594.900 4.000 596.820 4.280 ;
      LAYER met3 ;
        RECT 17.720 4.255 584.525 587.685 ;
      LAYER met4 ;
        RECT 214.585 61.375 250.050 420.745 ;
        RECT 252.450 61.375 253.350 420.745 ;
        RECT 255.750 61.375 256.650 420.745 ;
        RECT 259.050 61.375 259.950 420.745 ;
        RECT 262.350 61.375 326.850 420.745 ;
        RECT 329.250 61.375 330.150 420.745 ;
        RECT 332.550 61.375 333.450 420.745 ;
        RECT 335.850 61.375 336.750 420.745 ;
        RECT 339.150 61.375 403.650 420.745 ;
        RECT 406.050 61.375 406.950 420.745 ;
        RECT 409.350 61.375 410.250 420.745 ;
        RECT 412.650 61.375 413.550 420.745 ;
        RECT 415.950 61.375 433.875 420.745 ;
  END
END DSP48
END LIBRARY

