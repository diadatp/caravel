* NGSPICE file created from user_proj_example.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 D Q CLK VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 HI LO VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2oi_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2oi_4 A1_N A2_N B1 B2 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D X VGND VPWR
.ends

.subckt user_proj_example io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104]
+ la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109]
+ la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114]
+ la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119]
+ la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124]
+ la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69]
+ la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74]
+ la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7]
+ la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85]
+ la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90]
+ la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96]
+ la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10]
+ la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114]
+ la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119]
+ la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123]
+ la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57]
+ la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62]
+ la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67]
+ la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72]
+ la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77]
+ la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82]
+ la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87]
+ la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92]
+ la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97]
+ la_data_out[98] la_data_out[99] la_data_out[9] la_oen[0] la_oen[100] la_oen[101]
+ la_oen[102] la_oen[103] la_oen[104] la_oen[105] la_oen[106] la_oen[107] la_oen[108]
+ la_oen[109] la_oen[10] la_oen[110] la_oen[111] la_oen[112] la_oen[113] la_oen[114]
+ la_oen[115] la_oen[116] la_oen[117] la_oen[118] la_oen[119] la_oen[11] la_oen[120]
+ la_oen[121] la_oen[122] la_oen[123] la_oen[124] la_oen[125] la_oen[126] la_oen[127]
+ la_oen[12] la_oen[13] la_oen[14] la_oen[15] la_oen[16] la_oen[17] la_oen[18] la_oen[19]
+ la_oen[1] la_oen[20] la_oen[21] la_oen[22] la_oen[23] la_oen[24] la_oen[25] la_oen[26]
+ la_oen[27] la_oen[28] la_oen[29] la_oen[2] la_oen[30] la_oen[31] la_oen[32] la_oen[33]
+ la_oen[34] la_oen[35] la_oen[36] la_oen[37] la_oen[38] la_oen[39] la_oen[3] la_oen[40]
+ la_oen[41] la_oen[42] la_oen[43] la_oen[44] la_oen[45] la_oen[46] la_oen[47] la_oen[48]
+ la_oen[49] la_oen[4] la_oen[50] la_oen[51] la_oen[52] la_oen[53] la_oen[54] la_oen[55]
+ la_oen[56] la_oen[57] la_oen[58] la_oen[59] la_oen[5] la_oen[60] la_oen[61] la_oen[62]
+ la_oen[63] la_oen[64] la_oen[65] la_oen[66] la_oen[67] la_oen[68] la_oen[69] la_oen[6]
+ la_oen[70] la_oen[71] la_oen[72] la_oen[73] la_oen[74] la_oen[75] la_oen[76] la_oen[77]
+ la_oen[78] la_oen[79] la_oen[7] la_oen[80] la_oen[81] la_oen[82] la_oen[83] la_oen[84]
+ la_oen[85] la_oen[86] la_oen[87] la_oen[88] la_oen[89] la_oen[8] la_oen[90] la_oen[91]
+ la_oen[92] la_oen[93] la_oen[94] la_oen[95] la_oen[96] la_oen[97] la_oen[98] la_oen[99]
+ la_oen[9] wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12]
+ wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18]
+ wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23]
+ wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29]
+ wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5]
+ wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10]
+ wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16]
+ wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21]
+ wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27]
+ wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3]
+ wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0]
+ wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15]
+ wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20]
+ wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26]
+ wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31]
+ wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9]
+ wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i VPWR VGND
XFILLER_80_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_266 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_439 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_556 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_581 VGND VPWR sky130_fd_sc_hd__fill_1
X_6914_ _6866_/A _6865_/X _6914_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XPHY_3109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_601 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_1014 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_1134 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_623 VGND VPWR sky130_fd_sc_hd__decap_12
X_6845_ _6843_/Y _6844_/Y _6845_/X VGND VPWR sky130_fd_sc_hd__and2_4
XPHY_2419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1058 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_628 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_757 VGND VPWR sky130_fd_sc_hd__decap_12
X_6776_ _6770_/A _6769_/X _6776_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XPHY_1729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_959 VGND VPWR sky130_fd_sc_hd__decap_12
X_3988_ _7303_/A _3988_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_149_842 VGND VPWR sky130_fd_sc_hd__decap_12
X_5727_ _5696_/X _5699_/X _5700_/X _5727_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_148_385 VGND VPWR sky130_fd_sc_hd__decap_12
X_5658_ _5656_/X _5657_/X _5658_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_175_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1069 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1020 VGND VPWR sky130_fd_sc_hd__decap_12
X_4609_ _4609_/A _4565_/B _4609_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_190_141 VGND VPWR sky130_fd_sc_hd__decap_12
X_5589_ _5185_/A _4631_/B _5589_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_151_517 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_208 VGND VPWR sky130_fd_sc_hd__decap_12
X_7328_ io_in[17] _7329_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_117_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_411 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1143 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_455 VGND VPWR sky130_fd_sc_hd__decap_3
X_7259_ _7259_/A _7260_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_105_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_477 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_501 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_98 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1243 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1261 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_450 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_483 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_239 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_494 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_606 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_111 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1158 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_105 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_948 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_987 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_678 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_115 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_609 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_661 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_812 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_363 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_503 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_873 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_1024 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_867 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_664 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1008 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_1227 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_775 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_572 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_414 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_586 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_203 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_367 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_342 VGND VPWR sky130_fd_sc_hd__decap_12
X_4960_ _4958_/X _4959_/X _4958_/X _4959_/X _4960_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_149_1148 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_781 VGND VPWR sky130_fd_sc_hd__decap_12
X_3911_ _7321_/A _3911_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_205_562 VGND VPWR sky130_fd_sc_hd__decap_12
X_4891_ _4891_/A _4891_/B _4891_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_177_403 VGND VPWR sky130_fd_sc_hd__decap_12
X_6630_ _6630_/A _6630_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_3842_ _3842_/A _3843_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_60_795 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_626 VGND VPWR sky130_fd_sc_hd__decap_12
X_6561_ _6586_/A _6553_/X _6560_/Y _6561_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_3773_ _4512_/A _3773_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_201_790 VGND VPWR sky130_fd_sc_hd__decap_3
X_5512_ _5463_/X _5500_/X _5510_/X _5511_/X _5512_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_125_1192 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_171 VGND VPWR sky130_fd_sc_hd__decap_12
X_6492_ _7712_/Q _6492_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_146_845 VGND VPWR sky130_fd_sc_hd__decap_8
X_5443_ _4459_/A _5443_/B _5444_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_172_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_815 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_208 VGND VPWR sky130_fd_sc_hd__decap_12
X_5374_ _5359_/X _5365_/X _5372_/X _5373_/X _5374_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_7113_ _7628_/Q la_data_in[90] _7048_/X _7113_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_4325_ _4286_/X _4287_/X _4286_/X _4287_/X _4325_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_141_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_306 VGND VPWR sky130_fd_sc_hd__decap_12
X_7044_ la_data_in[91] _7044_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4256_ _4245_/X _4246_/X _4245_/X _4246_/X _4256_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_102_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_469 VGND VPWR sky130_fd_sc_hd__decap_12
X_4187_ _4171_/X _4174_/X _4187_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_110_970 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1174 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_910 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_386 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_39 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_239 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_701 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_965 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_521 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_464 VGND VPWR sky130_fd_sc_hd__decap_12
X_6828_ _7661_/Q _6830_/A VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_114 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6759_ _6736_/Y _6737_/Y _6758_/X _6759_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XPHY_1559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_525 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_461 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_995 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_848 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1030 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_1090 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_775 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_572 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_637 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1096 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_1260 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_607 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_1252 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_320 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_394 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_556 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_337 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_228 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_792 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_550 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_291 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_431 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_751 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1072 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1023 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_745 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1094 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_42_784 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_261 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1029 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_970 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_653 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_325 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_712 VGND VPWR sky130_fd_sc_hd__decap_12
X_4110_ _4092_/A _4091_/X _4092_/X _4110_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_151_1005 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_594 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_648 VGND VPWR sky130_fd_sc_hd__decap_12
X_5090_ _5077_/X _5083_/X _5077_/X _5083_/X _5090_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_190_1076 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_778 VGND VPWR sky130_fd_sc_hd__decap_12
X_4041_ _4010_/X _4011_/X _4010_/X _4011_/X _4041_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_84_618 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_383 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_164 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_175 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_876 VGND VPWR sky130_fd_sc_hd__decap_12
X_7800_ _7800_/D _3850_/A _7801_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_5992_ _6269_/A _5990_/X _5819_/X _5991_/Y _5993_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_64_375 VGND VPWR sky130_fd_sc_hd__decap_12
X_7731_ _7731_/D _7731_/Q _7797_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_197_509 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_239 VGND VPWR sky130_fd_sc_hd__decap_12
X_4943_ _4811_/X _4815_/X _4810_/X _4816_/X _4943_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_127_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_902 VGND VPWR sky130_fd_sc_hd__decap_12
X_7662_ _6893_/X _6825_/A _7658_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_71_1017 VGND VPWR sky130_fd_sc_hd__decap_12
X_4874_ _4838_/X _4873_/X _4838_/X _4873_/X _4874_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_60_581 VGND VPWR sky130_fd_sc_hd__decap_12
X_6613_ la_data_in[26] _6613_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_3825_ _6333_/A _3832_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_7593_ _7593_/HI la_data_out[120] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_165_417 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_1131 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_165_428 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_1208 VGND VPWR sky130_fd_sc_hd__decap_12
X_6544_ _6515_/A _6515_/B _6515_/X _6543_/X _6544_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_3756_ _5304_/A _5069_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_146_631 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_642 VGND VPWR sky130_fd_sc_hd__decap_12
X_6475_ _6431_/A _6431_/B _6475_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_106_506 VGND VPWR sky130_fd_sc_hd__decap_12
X_3687_ _6144_/A _6190_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_174_995 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_623 VGND VPWR sky130_fd_sc_hd__decap_12
X_5426_ _5095_/A _5300_/B _5428_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_161_645 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_859 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1102 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_509 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_902 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1233 VGND VPWR sky130_fd_sc_hd__decap_12
X_5357_ _5338_/X _5346_/X _5338_/X _5346_/X _5357_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_160_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1203 VGND VPWR sky130_fd_sc_hd__decap_12
X_4308_ _4308_/A _4309_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_173_1274 VGND VPWR sky130_fd_sc_hd__decap_3
X_5288_ _5228_/X _5285_/X _5286_/X _5287_/X _5332_/A VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_141_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1179 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_147 VGND VPWR sky130_fd_sc_hd__decap_12
X_7027_ _7636_/Q la_data_in[66] _6964_/X _7027_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_4239_ _4237_/X _4238_/X _4236_/X _4239_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_87_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_353 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_684 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_312 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_509 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_323 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_44 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1089 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_879 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_902 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_520 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_389 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1267 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_929 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_373 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_53 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_990 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1013 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1024 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_995 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_483 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1125 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1057 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_954 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_550 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_412 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_72 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_821 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_35 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1066 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1137 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_356 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_520 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_863 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_261 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_581 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_55 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_373 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_586 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_776 VGND VPWR sky130_fd_sc_hd__decap_6
X_4590_ _4590_/A _4590_/B _4592_/A VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_1890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_973 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_961 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_770 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_461 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1089 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_471 VGND VPWR sky130_fd_sc_hd__decap_12
X_6260_ _5993_/D _5766_/X _5765_/A _6260_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_192_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_336 VGND VPWR sky130_fd_sc_hd__decap_8
X_5211_ _5153_/X _5210_/X _5153_/X _5210_/X _5211_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_157_1269 VGND VPWR sky130_fd_sc_hd__decap_8
X_6191_ _4814_/A _6117_/X _6190_/X _6191_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_142_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_328 VGND VPWR sky130_fd_sc_hd__decap_8
X_5142_ _5137_/X _5141_/X _5140_/X _5142_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_111_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1046 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1068 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_916 VGND VPWR sky130_fd_sc_hd__decap_12
X_5073_ _5234_/A _4641_/B _5073_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_69_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_586 VGND VPWR sky130_fd_sc_hd__decap_8
X_4024_ _4005_/X _4023_/X _4005_/X _4023_/X _4024_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_84_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_971 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1204 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_898 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_684 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_306 VGND VPWR sky130_fd_sc_hd__decap_12
X_5975_ _5974_/A _5973_/X _5974_/X _5975_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_80_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_507 VGND VPWR sky130_fd_sc_hd__decap_12
X_4926_ _4926_/A _4926_/B _4926_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7714_ _7714_/D _7714_/Q _7785_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_178_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_929 VGND VPWR sky130_fd_sc_hd__decap_8
X_4857_ _4857_/A _4856_/X _4857_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7645_ _7004_/X _7645_/Q _7754_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_178_575 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_501 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_231 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_765 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_776 VGND VPWR sky130_fd_sc_hd__decap_12
X_3808_ wbs_dat_i[12] _3822_/B _3808_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_7576_ _7576_/HI la_data_out[103] VGND VPWR sky130_fd_sc_hd__conb_1
X_4788_ _4786_/X _4787_/X _4786_/X _4787_/X _4788_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_197_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_269 VGND VPWR sky130_fd_sc_hd__decap_12
X_6527_ _6527_/A _6526_/Y _6527_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_119_664 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_141 VGND VPWR sky130_fd_sc_hd__decap_12
X_3739_ _3738_/X _3712_/X _3741_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_107_826 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1257 VGND VPWR sky130_fd_sc_hd__decap_12
X_6458_ _7725_/Q la_data_in[123] _6393_/X _6458_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_84_1219 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_27 VGND VPWR sky130_fd_sc_hd__decap_12
X_5409_ _5341_/A _4854_/B _5409_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_161_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_306 VGND VPWR sky130_fd_sc_hd__decap_12
X_6389_ la_data_in[124] _6390_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_0_614 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_102_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1074 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_862 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_776 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_810 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_1088 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1214 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_662 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_301 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_98 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1072 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_63 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_581 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_703 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_726 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_586 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1067 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_242 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_776 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1168 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_224 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_567 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_297 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_973 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_73 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_721 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_391 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_1185 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_908 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_802 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_824 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_312 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_654 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_985 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_687 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_518 VGND VPWR sky130_fd_sc_hd__fill_1
X_5760_ _5745_/X _5755_/X _5753_/X _5756_/X _5760_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_188_851 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_581 VGND VPWR sky130_fd_sc_hd__decap_12
X_4711_ _4587_/X _4710_/X _4587_/X _4710_/X _4711_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_5691_ _4678_/A _4491_/A _5691_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_175_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1178 VGND VPWR sky130_fd_sc_hd__decap_12
X_7430_ io_oeb[25] _7430_/LO VGND VPWR sky130_fd_sc_hd__conb_1
X_4642_ _4642_/A _4642_/B _4642_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_175_578 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_269 VGND VPWR sky130_fd_sc_hd__decap_12
X_7361_ _5058_/A _7349_/X _7360_/Y _7387_/A _7361_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_163_729 VGND VPWR sky130_fd_sc_hd__decap_3
X_4573_ _4568_/X _4572_/X _4568_/X _4572_/X _4573_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_128_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_623 VGND VPWR sky130_fd_sc_hd__decap_12
X_6312_ _6308_/X _6311_/X _6057_/A _6312_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_162_239 VGND VPWR sky130_fd_sc_hd__decap_12
X_7292_ _7783_/Q _7292_/B _7292_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_200_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_954 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_645 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1033 VGND VPWR sky130_fd_sc_hd__decap_4
X_6243_ _6197_/X _6198_/B _6197_/X _6198_/B _6243_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_144_998 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_829 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_306 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_19 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_220 VGND VPWR sky130_fd_sc_hd__decap_12
X_6174_ _4989_/X _6174_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_97_562 VGND VPWR sky130_fd_sc_hd__decap_12
X_5125_ _5125_/A _5125_/B _5125_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_57_404 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_724 VGND VPWR sky130_fd_sc_hd__decap_8
X_5056_ _4552_/A _4782_/B _5056_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_211_1241 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_960 VGND VPWR sky130_fd_sc_hd__decap_12
X_4007_ _3738_/A _3950_/B _4007_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_77_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_604 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_857 VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_1_0_1_wb_clk_i clkbuf_1_0_1_wb_clk_i/A clkbuf_1_0_1_wb_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_129_1135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_367 VGND VPWR sky130_fd_sc_hd__decap_12
X_5958_ _5186_/A _4532_/A _5957_/Y _5958_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_197_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_337 VGND VPWR sky130_fd_sc_hd__decap_12
X_4909_ _4907_/X _4908_/X _4907_/X _4908_/X _4909_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_178_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_5889_ _5887_/X _5888_/X _5889_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_187_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_562 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_534 VGND VPWR sky130_fd_sc_hd__decap_12
X_7628_ _7116_/X _7628_/Q _7729_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_194_854 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_595 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1040 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_601 VGND VPWR sky130_fd_sc_hd__decap_8
X_7559_ _7559_/HI la_data_out[86] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_88_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1133 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_689 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_840 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_916 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_466 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_895 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1022 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_632 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1099 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_637 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_676 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_175 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_849 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_326 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_340 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_351 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_362 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_373 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_384 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_395 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_83 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1151 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_577 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_239 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_5 _4505_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_773 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_261 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_648 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1050 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_702 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1094 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_757 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_779 VGND VPWR sky130_fd_sc_hd__decap_12
X_6930_ la_data_in[77] _6931_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_54_429 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_481 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_963 VGND VPWR sky130_fd_sc_hd__decap_12
X_6861_ _6858_/Y _6859_/Y _6858_/Y _6859_/Y _6861_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_5812_ _5809_/X _5811_/X _5809_/X _5811_/X _5812_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_22_315 VGND VPWR sky130_fd_sc_hd__decap_12
X_6792_ _6792_/A _6763_/X _6792_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_179_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_495 VGND VPWR sky130_fd_sc_hd__decap_12
X_5743_ _5729_/X _5735_/X _5729_/X _5735_/X _5743_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_194_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1073 VGND VPWR sky130_fd_sc_hd__decap_8
X_5674_ _5665_/X _5672_/X _5665_/X _5672_/X _5674_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_148_556 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_876 VGND VPWR sky130_fd_sc_hd__decap_8
X_4625_ _4625_/A _4625_/B _4628_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_7413_ io_oeb[8] _7413_/LO VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_163_515 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1098 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_846 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_1008 VGND VPWR sky130_fd_sc_hd__decap_8
X_7344_ io_in[20] _7345_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_4556_ _4553_/X _4554_/X _4555_/X _4556_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_191_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_762 VGND VPWR sky130_fd_sc_hd__fill_1
X_7275_ io_in[8] _7275_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_1_208 VGND VPWR sky130_fd_sc_hd__decap_8
X_4487_ _4486_/A _4485_/X _4530_/A _4495_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_1_219 VGND VPWR sky130_fd_sc_hd__decap_8
X_6226_ _6223_/Y _6225_/Y _5396_/Y _6228_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_132_968 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_871 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1191 VGND VPWR sky130_fd_sc_hd__decap_6
X_6157_ _5032_/A _6155_/X _6101_/X _6157_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_106_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1172 VGND VPWR sky130_fd_sc_hd__decap_3
X_5108_ _3813_/X _4497_/B _5108_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_131_1036 VGND VPWR sky130_fd_sc_hd__fill_1
X_6088_ _6311_/B _6219_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_5039_ _5039_/A _6019_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_100_898 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_930 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_56 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_654 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_805 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_602 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_917 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_849 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_635 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_43 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1151 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1113 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_692 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1015 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_910 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_86 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_879 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_764 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_618 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_798 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1253 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1144 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_587 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_738 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_607 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_955 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1076 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1027 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_977 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_819 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_93 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_170 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_178 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_192 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_865 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_864 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_397 VGND VPWR sky130_fd_sc_hd__decap_12
X_4410_ _3738_/A _4459_/B _4410_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_8_396 VGND VPWR sky130_fd_sc_hd__fill_1
X_5390_ _5336_/X _5380_/X _5336_/X _5380_/X _5390_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_173_879 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_740 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_507 VGND VPWR sky130_fd_sc_hd__decap_12
X_4341_ _4327_/X _4333_/X _4339_/X _4340_/X _4341_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_158_1183 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_1134 VGND VPWR sky130_fd_sc_hd__fill_2
X_7060_ _7058_/Y _7060_/B _7060_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_4272_ _4270_/X _4271_/X _4270_/X _4271_/X _4272_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_1088 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_819 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1099 VGND VPWR sky130_fd_sc_hd__decap_12
X_6011_ _5547_/Y _6011_/B _6004_/Y _6010_/Y _6011_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_154_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_489 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_278 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_6913_ _6913_/A _6923_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_82_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_440 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1146 VGND VPWR sky130_fd_sc_hd__decap_12
X_6844_ la_data_in[54] _6844_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_51_944 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_714 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_202 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_938 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1029 VGND VPWR sky130_fd_sc_hd__decap_8
X_3987_ _3985_/Y _3986_/Y _3985_/Y _3986_/Y _3987_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6775_ _6885_/A _6773_/Y _6775_/C _6775_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_211_769 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_307 VGND VPWR sky130_fd_sc_hd__decap_12
X_5726_ _5715_/X _5716_/X _5715_/X _5716_/X _5726_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_148_331 VGND VPWR sky130_fd_sc_hd__decap_4
X_5657_ _5645_/X _5646_/X _5647_/X _5657_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_108_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1032 VGND VPWR sky130_fd_sc_hd__decap_4
X_4608_ _4605_/X _4606_/X _4813_/A _4608_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_5588_ _5585_/X _5586_/X _5587_/X _5588_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_163_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1111 VGND VPWR sky130_fd_sc_hd__decap_12
X_4539_ _4539_/A _4793_/B _4539_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7327_ _7327_/A _7321_/B _7327_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_104_423 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1155 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1245 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_220 VGND VPWR sky130_fd_sc_hd__decap_12
X_7258_ _7258_/A _7253_/B _7259_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_77_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_318 VGND VPWR sky130_fd_sc_hd__decap_12
X_6209_ _5565_/X _6201_/B _6209_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_104_489 VGND VPWR sky130_fd_sc_hd__decap_3
X_7189_ _7237_/A _7237_/B _7238_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_58_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_373 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_727 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_524 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1161 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_1233 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_952 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_708 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_440 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1273 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_4367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1246 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_281 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1268 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_123 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1227 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_117 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_999 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_178 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_257 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_52 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_802 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_824 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_375 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_812 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_805 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1036 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1058 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1203 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_550 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_787 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_638 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_521 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_841 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_448 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_220 VGND VPWR sky130_fd_sc_hd__decap_12
X_3910_ _7343_/A _3910_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_32_410 VGND VPWR sky130_fd_sc_hd__decap_12
X_4890_ _4885_/X _4889_/X _4885_/X _4889_/X _4891_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_205_574 VGND VPWR sky130_fd_sc_hd__decap_12
X_3841_ _3832_/A _3841_/B _3840_/Y _7802_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_177_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_977 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_638 VGND VPWR sky130_fd_sc_hd__decap_3
X_3772_ _4844_/A _4512_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_6560_ _6560_/A _6553_/B _6560_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_125_1160 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_971 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_802 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_418 VGND VPWR sky130_fd_sc_hd__fill_2
X_5511_ _5463_/X _5500_/X _5463_/X _5500_/X _5511_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_192_429 VGND VPWR sky130_fd_sc_hd__decap_12
X_6491_ _6190_/A _6885_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_9_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1106 VGND VPWR sky130_fd_sc_hd__decap_8
X_5442_ _5442_/A _5442_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_145_367 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_529 VGND VPWR sky130_fd_sc_hd__decap_12
X_5373_ _5359_/X _5365_/X _5359_/X _5365_/X _5373_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_126_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_337 VGND VPWR sky130_fd_sc_hd__decap_12
X_4324_ _4305_/X _4306_/X _4305_/X _4306_/X _4324_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7112_ _7091_/X _7110_/X _7111_/Y _7629_/D VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_113_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_540 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_318 VGND VPWR sky130_fd_sc_hd__decap_8
X_7043_ _7043_/A _7043_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4255_ _4248_/Y _4249_/X _4248_/Y _4249_/X _4255_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_87_638 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1120 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1014 VGND VPWR sky130_fd_sc_hd__decap_8
X_4186_ _4180_/X _4185_/X _4179_/X _4186_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_132_1142 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1025 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_982 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_513 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1186 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_226 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_398 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_410 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_916 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_977 VGND VPWR sky130_fd_sc_hd__decap_12
X_6827_ _6825_/Y _6827_/B _6827_/X VGND VPWR sky130_fd_sc_hd__and2_4
XPHY_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_476 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1230 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1121 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6758_ _6738_/X _6758_/B _6758_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_177_960 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_126 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_407 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1274 VGND VPWR sky130_fd_sc_hd__decap_3
X_5709_ _5709_/A _5709_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_164_610 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_6689_ _6624_/A la_data_in[22] _6626_/X _6689_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_12_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_473 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_826 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_325 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_754 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_871 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1053 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_787 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_144_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_735 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1272 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_705 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_502 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1256 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1215 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_373 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_30 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1237 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_877 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_568 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1052 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_404 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_977 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_903 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1035 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_62 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_544 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_448 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1049 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_947 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_802 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_982 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_620 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_665 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_925 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_724 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1017 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_381 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1088 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_12_0_wb_clk_i clkbuf_3_6_0_wb_clk_i/X _7801_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4040_ _4013_/X _4022_/X _4013_/X _4022_/X _4040_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_204_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_833 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_395 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_535 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_343 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_663 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_803 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_888 VGND VPWR sky130_fd_sc_hd__decap_12
X_5991_ _5820_/A _5856_/Y _5991_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_80_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_861 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_387 VGND VPWR sky130_fd_sc_hd__decap_3
X_7730_ _6381_/Y _7730_/Q _7801_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_91_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_398 VGND VPWR sky130_fd_sc_hd__fill_1
X_4942_ _4874_/X _4875_/X _4817_/X _4876_/X _4942_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_17_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1233 VGND VPWR sky130_fd_sc_hd__decap_12
X_7661_ _6896_/X _7661_/Q _7658_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_178_735 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_914 VGND VPWR sky130_fd_sc_hd__fill_1
X_4873_ _4871_/X _4872_/X _4871_/X _4872_/X _4873_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_251 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1029 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_413 VGND VPWR sky130_fd_sc_hd__decap_12
X_6612_ _6612_/A _6612_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_177_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_593 VGND VPWR sky130_fd_sc_hd__decap_12
X_3824_ _6144_/A _6333_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_159_960 VGND VPWR sky130_fd_sc_hd__fill_1
X_7592_ _7592_/HI la_data_out[119] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_192_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1143 VGND VPWR sky130_fd_sc_hd__decap_12
X_3755_ _4847_/A _5304_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_6543_ _6516_/Y _6518_/B _6518_/X _6542_/X _6543_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_146_654 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_440 VGND VPWR sky130_fd_sc_hd__decap_12
X_3686_ wb_rst_i _6144_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_6474_ _6432_/X _6472_/X _6473_/Y _6474_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_106_518 VGND VPWR sky130_fd_sc_hd__fill_1
X_5425_ _5420_/X _5424_/X _5423_/X _5425_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_161_635 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_161_657 VGND VPWR sky130_fd_sc_hd__decap_12
X_5356_ _5352_/X _5355_/X _5352_/X _5355_/X _5356_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_82_1114 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_807 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_829 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_1215 VGND VPWR sky130_fd_sc_hd__fill_1
X_4307_ _4257_/X _4288_/X _4305_/X _4306_/X _4307_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_88_947 VGND VPWR sky130_fd_sc_hd__decap_12
X_5287_ _5228_/X _5285_/X _5228_/X _5285_/X _5287_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_4238_ _4535_/A _4346_/B _4238_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7026_ _6971_/X _7023_/X _7025_/Y _7026_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_101_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_159 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_991 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_4169_ _4641_/B _4591_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_114_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_790 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_877 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_335 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_56 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_379 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1235 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_532 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_727 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_385 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_749 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_930 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1090 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1142 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_109_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1036 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1069 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_966 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_111 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_122 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_540 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_402 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_424 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_381 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_479 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1261 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_62 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_84 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1143 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1260 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_47 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1078 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1187 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_825 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1149 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_842 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_379 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_532 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_571 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_245 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_727 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_385 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_621 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1013 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_93 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_440 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_805 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_985 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_973 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_782 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_473 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_410 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_1264 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_2_1_wb_clk_i clkbuf_2_2_1_wb_clk_i/A clkbuf_2_2_1_wb_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_143_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1117 VGND VPWR sky130_fd_sc_hd__decap_12
X_5210_ _5195_/X _5209_/X _5195_/X _5209_/X _5210_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_143_668 VGND VPWR sky130_fd_sc_hd__decap_3
X_6190_ _6190_/A _6190_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_43_3 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_178 VGND VPWR sky130_fd_sc_hd__decap_12
X_5141_ _5140_/A _5140_/B _5140_/X _5141_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_124_893 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_733 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_532 VGND VPWR sky130_fd_sc_hd__decap_12
X_5072_ _5072_/A _4624_/B _5072_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_96_276 VGND VPWR sky130_fd_sc_hd__decap_6
X_4023_ _4006_/X _4012_/X _4013_/X _4022_/X _4023_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_96_298 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_844 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1216 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_471 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_324 VGND VPWR sky130_fd_sc_hd__decap_12
X_5974_ _5974_/A _5974_/B _5974_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_197_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_666 VGND VPWR sky130_fd_sc_hd__decap_6
X_7713_ _6558_/Y io_out[0] _7696_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4925_ _4553_/A _4925_/B _4926_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_100_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_532 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1041 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_733 VGND VPWR sky130_fd_sc_hd__decap_12
X_7644_ _7007_/X _7644_/Q _7754_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4856_ _4771_/A _4856_/B _4856_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_20_243 VGND VPWR sky130_fd_sc_hd__decap_12
X_3807_ _4589_/A _3798_/B _3807_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_21_788 VGND VPWR sky130_fd_sc_hd__decap_4
X_7575_ _7575_/HI la_data_out[102] VGND VPWR sky130_fd_sc_hd__conb_1
X_4787_ _4524_/X _4525_/X _4524_/X _4525_/X _4787_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_140_1252 VGND VPWR sky130_fd_sc_hd__decap_3
X_6526_ la_data_in[3] _6526_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_14_1266 VGND VPWR sky130_fd_sc_hd__decap_8
X_3738_ _3738_/A _3738_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_107_838 VGND VPWR sky130_fd_sc_hd__decap_12
X_6457_ _6440_/X _6454_/X _6456_/Y _6457_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_173_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_5408_ _5198_/A _4852_/B _5408_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_6388_ _7726_/Q _6390_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_161_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1050 VGND VPWR sky130_fd_sc_hd__decap_12
X_5339_ _5215_/A _4328_/B _5339_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_102_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_800 VGND VPWR sky130_fd_sc_hd__fill_1
X_7009_ _6923_/A _6981_/X _7008_/Y _7009_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_169_1108 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_611 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1002 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_830 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1141 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1084 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_75 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_812 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_593 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_715 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_215 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_788 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_236 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_259 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_41 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_771 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_985 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_85 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_410 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_679 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_508 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_965 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_616 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_987 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1209 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1197 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_928 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_373 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_901 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_129 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_8_1091 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_956 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_836 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_997 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_699 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_880 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1233 VGND VPWR sky130_fd_sc_hd__decap_12
X_4710_ _4691_/X _4709_/X _4691_/X _4709_/X _4710_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_188_863 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_593 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1263 VGND VPWR sky130_fd_sc_hd__decap_12
X_5690_ _5687_/X _5688_/X _5689_/X _5690_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_175_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1119 VGND VPWR sky130_fd_sc_hd__decap_8
X_4641_ _5130_/A _4641_/B _4642_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_4572_ _4569_/X _4570_/X _4571_/X _4572_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_7360_ io_in[23] _7360_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_6311_ _5974_/X _6311_/B _6311_/C _6311_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_143_421 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_635 VGND VPWR sky130_fd_sc_hd__decap_6
X_7291_ _7259_/A _7292_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_7_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_657 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_123 VGND VPWR sky130_fd_sc_hd__decap_12
X_6242_ _6240_/Y _6242_/B _6242_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_170_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_785 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_1253 VGND VPWR sky130_fd_sc_hd__decap_3
X_6173_ _6089_/X _6171_/X _6172_/X _6173_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_44_1215 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_232 VGND VPWR sky130_fd_sc_hd__decap_12
X_5124_ _4505_/A _4485_/B _5125_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_97_574 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_416 VGND VPWR sky130_fd_sc_hd__decap_8
X_5055_ _5052_/X _5053_/X _5054_/X _5055_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_211_1253 VGND VPWR sky130_fd_sc_hd__decap_12
X_4006_ _3976_/X _3977_/X _3976_/X _3977_/X _4006_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_66_972 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1013 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_825 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_616 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1008 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_986 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_379 VGND VPWR sky130_fd_sc_hd__decap_12
X_5957_ _7747_/Q _5957_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_209_1160 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_198 VGND VPWR sky130_fd_sc_hd__decap_12
X_4908_ _4828_/X _4832_/X _4831_/X _4908_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_194_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_349 VGND VPWR sky130_fd_sc_hd__decap_12
X_5888_ _5787_/A _4480_/Y _5888_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_178_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_7627_ _7118_/X _7627_/Q _7729_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4839_ _4631_/X _4635_/X _4634_/X _4839_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_166_546 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_866 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_440 VGND VPWR sky130_fd_sc_hd__decap_6
X_7558_ _7558_/HI la_data_out[85] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_119_462 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1120 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_1142 VGND VPWR sky130_fd_sc_hd__decap_12
X_6509_ _6507_/Y _6508_/Y _6507_/Y _6508_/Y _6575_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_140_1093 VGND VPWR sky130_fd_sc_hd__decap_12
X_7489_ _7489_/HI la_data_out[16] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_4_239 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1145 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1167 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_412 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_852 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_703 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_75 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1001 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_641 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1072 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_717 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1034 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_1094 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_975 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_666 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_688 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_330 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_891 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_341 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_352 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_363 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_374 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_385 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_642 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_396 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_62 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_596 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_95 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_760 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_1163 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_922 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_398 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_6 _4562_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_1204 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_251 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_785 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_773 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_349 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_511 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_438 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_1270 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_764 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_633 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_184 VGND VPWR sky130_fd_sc_hd__decap_12
X_6860_ _6860_/A la_data_in[48] _6922_/A VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_63_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1219 VGND VPWR sky130_fd_sc_hd__fill_1
X_5811_ _5801_/X _5810_/X _5801_/X _5810_/X _5811_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_614 VGND VPWR sky130_fd_sc_hd__decap_12
X_6791_ _6913_/A _6795_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_22_327 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_159 VGND VPWR sky130_fd_sc_hd__decap_12
X_5742_ _5739_/X _5740_/X _5749_/B _5742_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_176_800 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_872 VGND VPWR sky130_fd_sc_hd__fill_2
X_5673_ _5641_/X _5642_/X _5641_/X _5642_/X _5673_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_148_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_382 VGND VPWR sky130_fd_sc_hd__decap_12
X_7412_ io_oeb[7] _7412_/LO VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_124_1077 VGND VPWR sky130_fd_sc_hd__fill_2
X_4624_ _5052_/A _4624_/B _4624_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_50_1252 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_527 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1178 VGND VPWR sky130_fd_sc_hd__decap_12
X_7343_ _7343_/A _7321_/B _7343_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_144_730 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_421 VGND VPWR sky130_fd_sc_hd__decap_12
X_4555_ _4553_/X _4554_/X _4555_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_117_977 VGND VPWR sky130_fd_sc_hd__decap_12
X_7274_ _7780_/Q _7260_/B _7274_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_4486_ _4486_/A _4485_/X _4530_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_132_947 VGND VPWR sky130_fd_sc_hd__decap_8
X_6225_ _6225_/A _6225_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_103_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1072 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_703 VGND VPWR sky130_fd_sc_hd__decap_6
X_6156_ _5032_/A _6155_/X _6156_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_98_883 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_725 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_991 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1004 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1067 VGND VPWR sky130_fd_sc_hd__fill_1
X_5107_ _5099_/X _5103_/X _5099_/X _5103_/X _5107_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_44_1078 VGND VPWR sky130_fd_sc_hd__decap_12
X_6087_ _6087_/A _6087_/B _7787_/D VGND VPWR sky130_fd_sc_hd__nor2_4
X_5038_ _5027_/X _5028_/X _5027_/X _5028_/X _5040_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_57_279 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_419 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_227 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_791 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_942 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_68 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_666 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_452 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_817 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_3837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_11 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1172 VGND VPWR sky130_fd_sc_hd__decap_6
X_6989_ io_out[4] _6988_/X _6991_/B VGND VPWR sky130_fd_sc_hd__xnor2_4
XPHY_3859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_55 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_660 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_77 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_513 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1125 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1136 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1027 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1199 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_922 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_730 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_977 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_988 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_722 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_593 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_242 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_660 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1134 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_1265 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1156 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_235 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_514 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_964 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_666 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_435 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_468 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1088 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_1039 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_135 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_160 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_129 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_171 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_877 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_505 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_876 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_696 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_752 VGND VPWR sky130_fd_sc_hd__decap_8
X_4340_ _4327_/X _4333_/X _4327_/X _4333_/X _4340_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_1034 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_1056 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_581 VGND VPWR sky130_fd_sc_hd__decap_12
X_4271_ _4568_/A _4923_/B _4271_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_113_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1168 VGND VPWR sky130_fd_sc_hd__fill_2
X_6010_ _5584_/X _6010_/B _6010_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_140_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_330 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_419 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_780 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_227 VGND VPWR sky130_fd_sc_hd__decap_12
X_6912_ _6912_/A _6868_/X _6912_/C _6912_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_78_1130 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_452 VGND VPWR sky130_fd_sc_hd__decap_12
X_6843_ _6843_/A _6843_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_63_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_956 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_647 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_211_726 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1128 VGND VPWR sky130_fd_sc_hd__fill_1
X_6774_ la_data_in[47] _6774_/B _6775_/C VGND VPWR sky130_fd_sc_hd__and2_4
XPHY_1709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1188 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_669 VGND VPWR sky130_fd_sc_hd__fill_2
X_3986_ _3943_/X _3946_/Y _3958_/B _3986_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
X_5725_ _5718_/X _5719_/X _5718_/X _5719_/X _5725_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_10_319 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_855 VGND VPWR sky130_fd_sc_hd__decap_12
X_5656_ _5472_/X _5473_/X _5474_/X _5656_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_164_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_611 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_398 VGND VPWR sky130_fd_sc_hd__decap_12
X_4607_ _4605_/X _4606_/X _4813_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_5587_ _5585_/X _5586_/X _5587_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_50_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_154 VGND VPWR sky130_fd_sc_hd__decap_12
X_7326_ _5754_/A _7309_/X _7321_/X _7325_/Y wbs_dat_o[10] VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_163_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1123 VGND VPWR sky130_fd_sc_hd__decap_6
X_4538_ _4538_/A _4538_/B _4538_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_2_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_880 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_529 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_744 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_435 VGND VPWR sky130_fd_sc_hd__decap_12
X_7257_ _7388_/A _7257_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_89_135 VGND VPWR sky130_fd_sc_hd__decap_12
X_4469_ _4590_/A _4597_/B _4469_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_131_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_6208_ _6208_/A _6211_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_132_788 VGND VPWR sky130_fd_sc_hd__fill_1
X_7188_ _7175_/Y _7177_/B _7177_/X _7187_/X _7237_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_86_831 VGND VPWR sky130_fd_sc_hd__fill_1
X_6139_ _6139_/A _6319_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_85_330 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_652 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_566 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_886 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_739 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_536 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_791 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_4313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_711 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_964 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_32 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_733 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1233 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_4368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_945 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1258 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_956 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_619 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_276 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_129 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_269 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_86 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_471 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_155_836 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_696 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_482 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_313 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_387 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_508 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_809 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_606 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_991 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_536 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1199 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_271 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_731 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_422 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_967 VGND VPWR sky130_fd_sc_hd__decap_8
X_3840_ wbs_dat_i[8] _3848_/B _3840_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_38_1191 VGND VPWR sky130_fd_sc_hd__decap_3
X_3771_ _3771_/A _4844_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_34_1044 VGND VPWR sky130_fd_sc_hd__decap_12
X_5510_ _5505_/X _5509_/X _5505_/X _5509_/X _5510_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_814 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_983 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_190 VGND VPWR sky130_fd_sc_hd__decap_12
X_6490_ _6466_/X _6487_/A _6489_/X _7714_/D VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_158_685 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1036 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_184 VGND VPWR sky130_fd_sc_hd__decap_12
X_5441_ _5428_/X _5431_/X _5442_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_195_1137 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_1148 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_154 VGND VPWR sky130_fd_sc_hd__decap_12
X_5372_ _5371_/A _5370_/X _5371_/X _5372_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_7111_ _7091_/X _7110_/X _7024_/X _7111_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_126_593 VGND VPWR sky130_fd_sc_hd__decap_12
X_4323_ _4311_/Y _4312_/X _4311_/Y _4312_/X _4323_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_160_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_755 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_232 VGND VPWR sky130_fd_sc_hd__decap_12
X_7042_ _7040_/Y _7041_/Y _7042_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_141_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_788 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_4254_ _4251_/A _4250_/X _4447_/A _4316_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_80_1020 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_1004 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_330 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1184 VGND VPWR sky130_fd_sc_hd__decap_12
X_4185_ _4583_/A _4346_/B _4185_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_95_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_205 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_994 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_238 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_59 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_422 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6826_ la_data_in[60] _6827_/B VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_2229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_241 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_736 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_989 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1160 VGND VPWR sky130_fd_sc_hd__decap_12
X_6757_ _6739_/Y _6740_/Y _6756_/X _6758_/B VGND VPWR sky130_fd_sc_hd__o21a_4
XPHY_1539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_285 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1242 VGND VPWR sky130_fd_sc_hd__decap_12
X_3969_ _3913_/Y _3961_/X _3962_/X _3991_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_195_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_419 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_138 VGND VPWR sky130_fd_sc_hd__decap_12
X_5708_ _5602_/A _5443_/B _5709_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_52_1166 VGND VPWR sky130_fd_sc_hd__decap_12
X_6688_ _6651_/X _6686_/X _6687_/Y _7689_/D VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_176_482 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_56 VGND VPWR sky130_fd_sc_hd__decap_12
X_5639_ _5639_/A _5639_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_128_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_485 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_838 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_733 VGND VPWR sky130_fd_sc_hd__decap_8
X_7309_ _7256_/A _7309_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_160_883 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_831 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_747 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_514 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_818 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_42 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1249 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1064 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_4132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1097 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1017 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_74 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_769 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_589 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_814 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_994 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_825 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_953 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_632 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_560 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1080 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_175 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_937 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1029 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_370 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_393 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_447 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_381 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_392 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_845 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_547 VGND VPWR sky130_fd_sc_hd__fill_2
X_5990_ _5857_/X _5990_/B _5990_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_92_675 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_815 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_761 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1111 VGND VPWR sky130_fd_sc_hd__decap_12
X_4941_ _4892_/X _4940_/X _4892_/X _4940_/X _4941_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_206_873 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_293 VGND VPWR sky130_fd_sc_hd__decap_12
X_7660_ _7660_/D _7660_/Q _7658_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_162_1114 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1117 VGND VPWR sky130_fd_sc_hd__decap_12
X_4872_ _4662_/X _4673_/X _4638_/X _4674_/X _4872_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_60_550 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1245 VGND VPWR sky130_fd_sc_hd__decap_8
X_6611_ _6611_/A _6611_/B _6611_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_3823_ _3791_/A _3821_/X _3822_/Y _3823_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_7591_ _7591_/HI la_data_out[118] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_425 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_257 VGND VPWR sky130_fd_sc_hd__decap_12
X_6542_ _6519_/Y _6520_/Y _6541_/X _6542_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_3754_ _4519_/A _4847_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_192_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1155 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_836 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_858 VGND VPWR sky130_fd_sc_hd__decap_12
X_6473_ _6432_/X _6472_/X _6455_/X _6473_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_173_452 VGND VPWR sky130_fd_sc_hd__decap_12
X_5424_ _5421_/X _5422_/X _5423_/X _5424_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_127_891 VGND VPWR sky130_fd_sc_hd__decap_12
X_5355_ _5353_/X _5354_/X _5353_/X _5354_/X _5355_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_161_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_703 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1126 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_819 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_403 VGND VPWR sky130_fd_sc_hd__decap_12
X_4306_ _4257_/X _4288_/X _4257_/X _4288_/X _4306_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_88_937 VGND VPWR sky130_fd_sc_hd__decap_8
X_5286_ _5280_/X _5281_/X _5279_/X _5282_/X _5286_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_88_959 VGND VPWR sky130_fd_sc_hd__decap_12
X_7025_ _6971_/X _7023_/X _7024_/X _7025_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_4237_ _4236_/A _4236_/B _4236_/X _4237_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_75_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_812 VGND VPWR sky130_fd_sc_hd__decap_12
X_4168_ _4612_/A _4590_/B _4168_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_67_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_141 VGND VPWR sky130_fd_sc_hd__decap_12
X_4099_ _4038_/Y _4068_/X _4067_/X _4099_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_43_517 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_388 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_130_68 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1044 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_241 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_747 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_11 VGND VPWR sky130_fd_sc_hd__fill_1
X_6809_ _6745_/A la_data_in[34] _6747_/X _6809_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XPHY_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1247 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_544 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7789_ _6067_/X _7327_/A _7785_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_44 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_397 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_430 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_964 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1004 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_806 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_379 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_978 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_669 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_585 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_393 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_609 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_970 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1273 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1100 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_428 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_1013 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_480 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1272 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_1155 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_506 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_59 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1109 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_196 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_764 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_701 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_712 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_544 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_3294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_257 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_419 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_227 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_666 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_817 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_997 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1205 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_485 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_647 VGND VPWR sky130_fd_sc_hd__decap_6
X_5140_ _5140_/A _5140_/B _5140_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_69_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_436 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_544 VGND VPWR sky130_fd_sc_hd__decap_4
X_5071_ _5062_/Y _5070_/X _5062_/Y _5070_/X _5071_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_4022_ _4014_/X _4020_/X _4021_/X _4022_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_38_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_856 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_141 VGND VPWR sky130_fd_sc_hd__decap_12
X_5973_ _5973_/A _5973_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_7712_ _6561_/X _7712_/Q _7696_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4924_ _4505_/A _4399_/B _4926_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_178_511 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1080 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_7643_ _7009_/X _7643_/Q _7754_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_127_1053 VGND VPWR sky130_fd_sc_hd__decap_12
X_4855_ _4000_/A _4856_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_60_380 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1097 VGND VPWR sky130_fd_sc_hd__fill_1
X_3806_ _5099_/A _4589_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_7574_ _7574_/HI la_data_out[101] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_255 VGND VPWR sky130_fd_sc_hd__decap_12
X_4786_ _4762_/X _4763_/X _4761_/X _4764_/X _4786_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_6525_ _6525_/A _6527_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_3737_ _4612_/A _3738_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_146_441 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1109 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_997 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_154 VGND VPWR sky130_fd_sc_hd__decap_12
X_6456_ _6440_/X _6454_/X _6455_/X _6456_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_173_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_349 VGND VPWR sky130_fd_sc_hd__decap_12
X_5407_ _5402_/X _5406_/X _5405_/X _5407_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_133_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_850 VGND VPWR sky130_fd_sc_hd__decap_4
X_6387_ _6387_/A _6387_/B _6387_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_86_1081 VGND VPWR sky130_fd_sc_hd__decap_12
X_5338_ _5237_/X _5238_/X _5239_/X _5338_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_173_1062 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1182 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_544 VGND VPWR sky130_fd_sc_hd__decap_12
X_5269_ _5114_/X _5115_/X _5114_/X _5115_/X _5269_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_130_886 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_7008_ _7008_/A _7008_/B _7008_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_75_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_44 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_867 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_450 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_601 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_366 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_163 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1170 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_196 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_842 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1153 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1044 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1096 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_566 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1115 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_87 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1058 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_391 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_419 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1069 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_846 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_727 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_536 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_227 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_110 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_53 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_647 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_742 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_764 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_989 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_861 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_786 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_872 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_999 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_894 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_820 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_498 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_715 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_9 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1081 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_968 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_910 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_612 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_848 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_965 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_155 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_550 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_892 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_875 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_1215 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_520 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1275 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_886 VGND VPWR sky130_fd_sc_hd__decap_12
X_4640_ _4640_/A _4625_/B _4642_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_175_525 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_396 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_430 VGND VPWR sky130_fd_sc_hd__decap_12
X_4571_ _4569_/X _4570_/X _4571_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_190_506 VGND VPWR sky130_fd_sc_hd__decap_12
X_6310_ _5969_/X _6309_/Y _6311_/C VGND VPWR sky130_fd_sc_hd__or2_4
X_7290_ _7750_/Q _7280_/X _7286_/X _7289_/Y wbs_dat_o[4] VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_171_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_135 VGND VPWR sky130_fd_sc_hd__decap_12
X_6241_ _5059_/Y _6117_/X _6190_/X _6242_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_144_978 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_669 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_466 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1008 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_6172_ _5020_/Y _6158_/X _6144_/X _6172_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_83_1276 VGND VPWR sky130_fd_sc_hd__fill_1
X_5123_ _4499_/A _5123_/B _5125_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_112_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1210 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_428 VGND VPWR sky130_fd_sc_hd__decap_12
X_5054_ _5052_/X _5053_/X _5054_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_38_642 VGND VPWR sky130_fd_sc_hd__decap_12
X_4005_ _4005_/A _3981_/X _4005_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_211_1265 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_984 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1142 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1025 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_837 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1058 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_628 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_818 VGND VPWR sky130_fd_sc_hd__decap_12
X_5956_ _5946_/A _5945_/X _5946_/Y _5956_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_111_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_1150 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_998 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_842 VGND VPWR sky130_fd_sc_hd__decap_12
X_4907_ _4905_/X _4906_/X _4905_/X _4906_/X _4907_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_5887_ _5731_/A _4477_/A _5887_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_33_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_812 VGND VPWR sky130_fd_sc_hd__decap_12
X_4838_ _4818_/X _4837_/X _4818_/X _4837_/X _4838_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7626_ _7626_/D _7626_/Q _7729_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_178_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1020 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_558 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_878 VGND VPWR sky130_fd_sc_hd__decap_6
X_7557_ _7557_/HI la_data_out[84] VGND VPWR sky130_fd_sc_hd__conb_1
X_4769_ _4769_/A _4512_/B _4769_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_140_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_208 VGND VPWR sky130_fd_sc_hd__decap_12
X_6508_ la_data_in[9] _6508_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_119_474 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_794 VGND VPWR sky130_fd_sc_hd__decap_8
X_7488_ _7488_/HI la_data_out[15] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_134_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1154 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_56 VGND VPWR sky130_fd_sc_hd__decap_12
X_6439_ _6396_/A _6396_/B _6396_/X _6438_/X _6439_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_162_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_820 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_959 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_435 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_907 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1040 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_87 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_707 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_653 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1261 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_729 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_1118 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_921 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_995 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1079 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_965 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_807 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_987 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_369 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1139 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_306 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_320 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_331 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_342 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_339 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_520 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_353 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_531 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_364 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_672 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_375 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_374 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_300 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_386 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_397 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1142 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_934 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_7 _4782_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1216 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_753 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_561 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_785 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_564 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_428 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_973 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_623 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_122 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_196 VGND VPWR sky130_fd_sc_hd__decap_12
X_5810_ _5751_/Y _5752_/X _5751_/Y _5752_/X _5810_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_762 VGND VPWR sky130_fd_sc_hd__fill_1
X_6790_ _6765_/X _6788_/X _6789_/Y _7676_/D VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_34_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_626 VGND VPWR sky130_fd_sc_hd__decap_12
X_5741_ _5739_/X _5740_/X _5749_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_210_418 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1050 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_672 VGND VPWR sky130_fd_sc_hd__decap_12
X_5672_ _5668_/X _5669_/X _5670_/X _5671_/X _5672_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_187_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_361 VGND VPWR sky130_fd_sc_hd__decap_8
X_7411_ io_oeb[6] _7411_/LO VGND VPWR sky130_fd_sc_hd__conb_1
X_4623_ _4595_/X _4599_/X _4598_/X _4623_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_30_394 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_208 VGND VPWR sky130_fd_sc_hd__decap_12
X_7342_ _5503_/A _7388_/A _7338_/X _7341_/Y wbs_dat_o[13] VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_163_539 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_1275 VGND VPWR sky130_fd_sc_hd__fill_2
X_4554_ _4554_/A _4597_/B _4554_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_116_433 VGND VPWR sky130_fd_sc_hd__decap_12
X_7273_ _7747_/Q _7257_/X _7269_/X _7272_/Y wbs_dat_o[1] VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_171_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_764 VGND VPWR sky130_fd_sc_hd__fill_1
X_4485_ _4485_/A _4485_/B _4485_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_89_306 VGND VPWR sky130_fd_sc_hd__decap_12
X_6224_ _6197_/X _6000_/B _6008_/B _6225_/A VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_106_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_6155_ _6147_/Y _6154_/Y _5030_/Y _6155_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_112_661 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1084 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_895 VGND VPWR sky130_fd_sc_hd__decap_12
X_5106_ _5092_/X _5105_/X _5092_/X _5105_/X _5106_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_131_1016 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_737 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_171 VGND VPWR sky130_fd_sc_hd__decap_12
X_6086_ _3993_/A _6084_/X _6085_/X _6087_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_39_940 VGND VPWR sky130_fd_sc_hd__decap_12
X_5037_ _5033_/X _5034_/X _5035_/X _5036_/X _5039_/A VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_45_409 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_910 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_4506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_239 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_954 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_948 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_678 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_3838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_464 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_306 VGND VPWR sky130_fd_sc_hd__decap_12
X_6988_ _6926_/Y _6927_/Y _6994_/B _6988_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_94_1180 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_1191 VGND VPWR sky130_fd_sc_hd__decap_12
X_5939_ _5938_/A _5937_/X _5938_/X _5940_/B VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_179_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1044 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_300 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_709 VGND VPWR sky130_fd_sc_hd__fill_1
X_7609_ _7230_/X _7609_/Q _7729_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_142_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_934 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_444 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_797 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_745 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_840 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_672 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_276 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_1168 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_556 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_247 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_718 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1062 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_526 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_902 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_166 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_447 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_80 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_150 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_172 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_171 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_183 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_361 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_194 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_517 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_888 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_764 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_915 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1054 VGND VPWR sky130_fd_sc_hd__fill_1
X_4270_ _4269_/A _4268_/X _4269_/X _4270_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_141_745 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_436 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_1079 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_593 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_458 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_501 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_409 VGND VPWR sky130_fd_sc_hd__fill_1
X_6911_ _6911_/A _6867_/X _6912_/C VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_54_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_943 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_954 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_464 VGND VPWR sky130_fd_sc_hd__decap_12
X_6842_ _6840_/Y _6842_/B _6842_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_62_250 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_907 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_581 VGND VPWR sky130_fd_sc_hd__decap_12
X_6773_ la_data_in[47] _6774_/B _6773_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_51_968 VGND VPWR sky130_fd_sc_hd__decap_8
X_3985_ _3918_/X _3924_/X _3926_/X _3985_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_211_738 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1142 VGND VPWR sky130_fd_sc_hd__decap_12
X_5724_ _5677_/X _5722_/A _5723_/X _5724_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_176_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_867 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_804 VGND VPWR sky130_fd_sc_hd__decap_12
X_5655_ _5498_/X _5499_/X _5498_/X _5499_/X _5655_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_191 VGND VPWR sky130_fd_sc_hd__decap_12
X_4606_ _4561_/A _4562_/B _4606_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_164_859 VGND VPWR sky130_fd_sc_hd__decap_3
X_5586_ _5233_/A _4277_/A _5586_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_175_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_731 VGND VPWR sky130_fd_sc_hd__fill_1
X_7325_ _5602_/A _7322_/X _7324_/X _7325_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
X_4537_ _4529_/Y _4536_/X _4529_/Y _4536_/X _4537_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_190_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_561 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1252 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1105 VGND VPWR sky130_fd_sc_hd__decap_12
X_7256_ _7256_/A _7388_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_144_594 VGND VPWR sky130_fd_sc_hd__decap_8
X_4468_ _4461_/A _4596_/B _4470_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_104_447 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_147 VGND VPWR sky130_fd_sc_hd__decap_12
X_6207_ _6207_/A _6206_/X _7769_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_137_1269 VGND VPWR sky130_fd_sc_hd__decap_8
X_7187_ _7180_/A _7180_/B _7180_/X _7186_/X _7187_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_4399_ _4512_/A _4399_/B _4400_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_131_277 VGND VPWR sky130_fd_sc_hd__fill_1
X_6138_ _6138_/A _6137_/X _6138_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_100_642 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_556 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_664 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_578 VGND VPWR sky130_fd_sc_hd__fill_2
X_6069_ _6208_/A _6185_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_22_1130 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1213 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_39 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_548 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_723 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_44 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1215 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_4358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_570 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1128 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_968 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_288 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_32 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_489 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_1062 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_848 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_494 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_325 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_656 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_764 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_285 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_745 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_15 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_26 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_618 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_501 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1041 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1033 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1093 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_1112 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_578 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_729 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1107 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_743 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_294 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_428 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1170 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_787 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1181 VGND VPWR sky130_fd_sc_hd__decap_8
X_3770_ _7810_/Q _3771_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_160_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_692 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_782 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_506 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_995 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_837 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_697 VGND VPWR sky130_fd_sc_hd__decap_4
X_5440_ _5401_/X _5418_/X _5438_/X _5439_/X _5440_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_9_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1050 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_347 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_5371_ _5371_/A _5370_/X _5371_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_172_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_317 VGND VPWR sky130_fd_sc_hd__decap_12
X_7110_ _7043_/A la_data_in[91] _7045_/X _7110_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_4322_ _4321_/X _4322_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_5_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_767 VGND VPWR sky130_fd_sc_hd__decap_8
X_7041_ la_data_in[92] _7041_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4253_ _4253_/A _4447_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_99_489 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1100 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_428 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1032 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1043 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_832 VGND VPWR sky130_fd_sc_hd__decap_12
X_4184_ _4459_/B _4346_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_45_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_718 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_898 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_835 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_868 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_559 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_751 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_283 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_7_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A clkbuf_3_7_0_wb_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_6825_ _6825_/A _6825_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_253 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1150 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_489 VGND VPWR sky130_fd_sc_hd__decap_12
X_3968_ _3993_/A _3962_/X _3968_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_6756_ _6741_/X _6804_/B _6756_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_91_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_297 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1254 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_269 VGND VPWR sky130_fd_sc_hd__decap_12
X_5707_ _5707_/A _5707_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_148_141 VGND VPWR sky130_fd_sc_hd__decap_12
X_6687_ _6651_/X _6686_/X _6670_/X _6687_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_192_910 VGND VPWR sky130_fd_sc_hd__decap_12
X_3899_ _3866_/X _3899_/B _3899_/C _7795_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_177_995 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_539 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_494 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1268 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1208 VGND VPWR sky130_fd_sc_hd__decap_12
X_5638_ _3813_/X _4793_/B _5638_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_12_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_807 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_806 VGND VPWR sky130_fd_sc_hd__fill_1
X_5569_ _5291_/X _5296_/X _5290_/X _5297_/X _5569_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_151_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_305 VGND VPWR sky130_fd_sc_hd__decap_4
X_7308_ _7753_/Q _7280_/X _7303_/X _7307_/Y wbs_dat_o[7] VGND VPWR sky130_fd_sc_hd__a211o_4
X_7239_ _7605_/Q la_data_in[99] _7177_/X _7239_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_144_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1088 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1222 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_759 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_331 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_662 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_802 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_718 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_312 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_54 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_239 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_98 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_531 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1087 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_581 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1029 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_776 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_86 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_962 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_1234 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_86 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_651 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_818 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_509 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_666 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_475 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1130 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_572 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1092 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1016 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_862 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1027 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_850 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_861 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_949 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_872 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_802 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_504 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_684 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_654 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_507 VGND VPWR sky130_fd_sc_hd__decap_12
X_4940_ _4938_/X _4939_/X _4938_/X _4939_/X _4940_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_80_849 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1123 VGND VPWR sky130_fd_sc_hd__decap_12
X_4871_ _4850_/X _4870_/X _4850_/X _4870_/X _4871_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_75_1167 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1126 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_776 VGND VPWR sky130_fd_sc_hd__decap_12
X_3822_ wbs_dat_i[10] _3822_/B _3822_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_6610_ la_data_in[27] _6611_/B VGND VPWR sky130_fd_sc_hd__inv_8
X_7590_ _7590_/HI la_data_out[117] VGND VPWR sky130_fd_sc_hd__conb_1
X_6541_ _6521_/X _6541_/B _6541_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_177_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_804 VGND VPWR sky130_fd_sc_hd__decap_12
X_3753_ _4614_/A _4519_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_20_459 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_239 VGND VPWR sky130_fd_sc_hd__decap_12
X_6472_ _7720_/Q la_data_in[118] _6408_/X _6472_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_5423_ _5421_/X _5422_/X _5423_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_161_604 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1252 VGND VPWR sky130_fd_sc_hd__decap_12
X_5354_ _5240_/X _5244_/X _5240_/X _5244_/X _5354_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1233 VGND VPWR sky130_fd_sc_hd__decap_12
X_4305_ _4301_/X _4302_/X _4304_/Y _4305_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_142_873 VGND VPWR sky130_fd_sc_hd__decap_12
X_5285_ _5229_/X _5273_/X _5283_/X _5284_/X _5285_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_173_1266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_726 VGND VPWR sky130_fd_sc_hd__decap_12
X_7024_ _6905_/A _7024_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4236_ _4236_/A _4236_/B _4236_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_4_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_269 VGND VPWR sky130_fd_sc_hd__decap_12
X_4167_ _4625_/B _4590_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_68_684 VGND VPWR sky130_fd_sc_hd__decap_12
X_4098_ _4029_/Y _4030_/X _4029_/Y _4030_/X _4098_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_55_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_507 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_529 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_581 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_337 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1245 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_776 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6808_ _6754_/X _6806_/X _6807_/Y _6808_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XPHY_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_759 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1078 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_354 VGND VPWR sky130_fd_sc_hd__decap_12
X_7788_ _6075_/Y _7321_/A _7746_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_426 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_567 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1062 VGND VPWR sky130_fd_sc_hd__decap_12
X_6739_ _7670_/Q _6739_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_165_910 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_461 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_656 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_1076 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_818 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1038 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_614 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_157 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_179 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_459 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_556 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1044 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_781 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1025 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1167 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_378 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_518 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_242 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_776 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_855 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_724 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_80 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_269 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_910 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_398 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_960 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_291 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_965 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_902 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1217 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_957 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_467 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1005 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1038 VGND VPWR sky130_fd_sc_hd__decap_8
X_5070_ _5068_/X _5069_/X _5068_/X _5069_/X _5070_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_81_1160 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_971 VGND VPWR sky130_fd_sc_hd__decap_12
X_4021_ _4014_/X _4020_/X _4021_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_77_481 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_172 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_868 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_518 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_996 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_389 VGND VPWR sky130_fd_sc_hd__decap_12
X_5972_ _5972_/A _5972_/B _5973_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_52_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_581 VGND VPWR sky130_fd_sc_hd__decap_12
X_7711_ _6564_/X _6495_/A _7707_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4923_ _3773_/X _4923_/B _4923_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_33_540 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_871 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1092 VGND VPWR sky130_fd_sc_hd__decap_12
X_7642_ _7012_/X _7642_/Q _7754_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4854_ _4514_/A _4854_/B _4857_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_127_1065 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_392 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_757 VGND VPWR sky130_fd_sc_hd__decap_8
X_3805_ _4461_/A _5099_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_4785_ _4768_/X _4774_/X _4783_/X _4784_/X _4785_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_7573_ _7573_/HI la_data_out[100] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_159_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_548 VGND VPWR sky130_fd_sc_hd__fill_1
X_3736_ _4479_/A _4612_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_6524_ _6522_/Y _6523_/Y _6522_/Y _6523_/Y _6524_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_101_1205 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_453 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_818 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_166 VGND VPWR sky130_fd_sc_hd__decap_12
X_6455_ _6190_/A _6455_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_109_59 VGND VPWR sky130_fd_sc_hd__fill_2
X_5406_ _5405_/A _5404_/X _5405_/X _5406_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_6386_ la_data_in[125] _6387_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_133_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1030 VGND VPWR sky130_fd_sc_hd__decap_6
X_5337_ _5249_/X _5250_/X _5249_/X _5250_/X _5337_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_161_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1161 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_1074 VGND VPWR sky130_fd_sc_hd__decap_12
X_5268_ _5246_/X _5247_/X _5245_/X _5248_/X _5268_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_87_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1099 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_556 VGND VPWR sky130_fd_sc_hd__decap_12
X_4219_ _4219_/A _4219_/B _4219_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7007_ _6982_/X _7005_/X _7006_/Y _7007_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_5199_ _5186_/A _3930_/A _5199_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_84_930 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_654 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_462 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1160 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_175 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1182 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_11 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_501 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1105 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_735 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_825 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1127 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_578 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_245 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_858 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_739 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_216 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_548 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_239 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_954 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_604 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_626 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_497 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_754 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_1250 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_798 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_489 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_1106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1070 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1104 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_167 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_898 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_537 VGND VPWR sky130_fd_sc_hd__decap_12
X_4570_ _4570_/A _4570_/B _4570_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_128_442 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_518 VGND VPWR sky130_fd_sc_hd__fill_1
X_6240_ _6240_/A _6240_/B _6240_/C _6240_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_115_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1096 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_478 VGND VPWR sky130_fd_sc_hd__decap_8
X_6171_ _5048_/X _6152_/X _5048_/X _6152_/X _6171_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_83_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1203 VGND VPWR sky130_fd_sc_hd__decap_12
X_5122_ _4503_/A _4493_/X _5122_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_112_865 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_109 VGND VPWR sky130_fd_sc_hd__decap_12
X_5053_ _5128_/A _4898_/D _5053_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_112_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1222 VGND VPWR sky130_fd_sc_hd__decap_12
X_4004_ _4189_/A _4123_/B _4005_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_38_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_996 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_27 VGND VPWR sky130_fd_sc_hd__decap_12
X_5955_ _5947_/X _5948_/X _5947_/X _5948_/X _5955_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_40_307 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1215 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_178 VGND VPWR sky130_fd_sc_hd__decap_12
X_4906_ _4565_/A _4906_/B _4906_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_5886_ _5872_/X _5873_/X _5874_/X _5886_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_7625_ _7123_/X _7055_/A _7624_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4837_ _4819_/X _4836_/X _4819_/X _4836_/X _4837_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_239 VGND VPWR sky130_fd_sc_hd__decap_12
X_7556_ _7556_/HI la_data_out[83] VGND VPWR sky130_fd_sc_hd__conb_1
X_4768_ _4512_/X _4516_/X _4512_/X _4516_/X _4768_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_101_1002 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1062 VGND VPWR sky130_fd_sc_hd__decap_6
X_6507_ _6507_/A _6507_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_3719_ _4821_/A _3720_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_119_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_626 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1035 VGND VPWR sky130_fd_sc_hd__fill_2
X_4699_ _4698_/A _4698_/B _4698_/X _4699_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_7487_ _7487_/HI la_data_out[14] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_161_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1177 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1008 VGND VPWR sky130_fd_sc_hd__decap_12
X_6438_ _6397_/Y _6398_/Y _6465_/B _6438_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_20_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_776 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_926 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_68 VGND VPWR sky130_fd_sc_hd__decap_12
X_6369_ _6190_/A _6381_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_1_937 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_832 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_948 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_738 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1052 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_665 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_1273 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_1047 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_607 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_819 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_999 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_310 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_98 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_318 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_321 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_332 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_370 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_343 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_354 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_365 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_543 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_684 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_376 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_387 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_386 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_312 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_398 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_740 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_8 _5275_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_979 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_573 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_595 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_797 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_274 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1020 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_576 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1231 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_719 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_131 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_755 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_977 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_668 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_134 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_808 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_178 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_638 VGND VPWR sky130_fd_sc_hd__decap_3
X_5740_ _4749_/A _4491_/A _5740_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_76_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1073 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1024 VGND VPWR sky130_fd_sc_hd__decap_8
X_5671_ _5629_/X _5630_/X _5629_/X _5630_/X _5671_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_175_312 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_1035 VGND VPWR sky130_fd_sc_hd__decap_12
X_7410_ io_oeb[5] _7410_/LO VGND VPWR sky130_fd_sc_hd__conb_1
X_4622_ _4588_/X _4621_/X _4588_/X _4621_/X _4622_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_175_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1081 VGND VPWR sky130_fd_sc_hd__decap_12
X_4553_ _4553_/A _4596_/B _4553_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7341_ _4467_/A _7322_/X _7340_/X _7341_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_156_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_445 VGND VPWR sky130_fd_sc_hd__decap_12
X_4484_ _4562_/B _4485_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_7272_ _5216_/A _7262_/X _7271_/X _7272_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_171_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_787 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_318 VGND VPWR sky130_fd_sc_hd__decap_12
X_6223_ _6223_/A _6223_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_106_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_6154_ _6153_/X _6154_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_174_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_673 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1096 VGND VPWR sky130_fd_sc_hd__fill_2
X_5105_ _5098_/X _5104_/X _5098_/X _5104_/X _5105_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6085_ _6068_/A _6085_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_131_1028 VGND VPWR sky130_fd_sc_hd__decap_8
X_5036_ _5033_/X _5034_/X _5033_/X _5034_/X _5036_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_39_952 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_730 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_4529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_281 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_966 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1141 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_3839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6987_ _6993_/A _6986_/X _6994_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_80_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_909 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_459 VGND VPWR sky130_fd_sc_hd__decap_12
X_5938_ _5938_/A _5937_/X _5938_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_22_852 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_684 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_931 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1056 VGND VPWR sky130_fd_sc_hd__decap_12
X_5869_ _5865_/X _5866_/X _5867_/Y _5868_/X _5869_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_139_537 VGND VPWR sky130_fd_sc_hd__decap_12
X_7608_ _7233_/X _7608_/Q _7729_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_194_654 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_816 VGND VPWR sky130_fd_sc_hd__decap_8
X_7539_ _7539_/HI la_data_out[66] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_182_849 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_990 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1250 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_852 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_1245 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_215 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_259 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_911 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_602 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_1074 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_538 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_292 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_947 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_1068 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_140 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_971 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_151 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_993 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_162 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_173 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_300 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_184 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_344 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_721 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1120 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1011 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1142 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_562 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_787 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_927 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1126 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_415 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_9_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/A _7797_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_207_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_297 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_822 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_833 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_911 VGND VPWR sky130_fd_sc_hd__decap_12
X_6910_ _6869_/X _6908_/X _6909_/Y _6910_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_94_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_281 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_966 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_903 VGND VPWR sky130_fd_sc_hd__decap_12
X_6841_ la_data_in[55] _6842_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_165_1135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1146 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_919 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_593 VGND VPWR sky130_fd_sc_hd__decap_8
X_6772_ io_out[2] _6771_/X _6774_/B VGND VPWR sky130_fd_sc_hd__xnor2_4
X_3984_ _3997_/A _3956_/X _3984_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_5723_ _5721_/Y _5722_/Y _5723_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_206_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_654 VGND VPWR sky130_fd_sc_hd__decap_6
X_5654_ _5644_/X _5653_/X _5644_/X _5653_/X _5654_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_164_816 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_676 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1160 VGND VPWR sky130_fd_sc_hd__decap_8
X_4605_ _3720_/A _5300_/B _4605_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_191_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1130 VGND VPWR sky130_fd_sc_hd__decap_12
X_5585_ _5341_/A _4145_/A _5585_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7324_ _7323_/Y _7324_/B _7324_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4536_ _4530_/X _4535_/X _4530_/X _4535_/X _4536_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_117_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_916 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_573 VGND VPWR sky130_fd_sc_hd__decap_6
X_7255_ _7354_/A _7256_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_176_1275 VGND VPWR sky130_fd_sc_hd__fill_2
X_4467_ _4467_/A _4595_/B _4467_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_172_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_59 VGND VPWR sky130_fd_sc_hd__fill_2
X_6206_ _4529_/Y _6117_/X _6190_/X _6206_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_131_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_459 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_159 VGND VPWR sky130_fd_sc_hd__decap_12
X_4398_ _4769_/A _4925_/B _4400_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_7186_ _7181_/Y _7182_/Y _7246_/B _7186_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_6137_ _6024_/Y _4451_/X _4443_/X _6137_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_112_492 VGND VPWR sky130_fd_sc_hd__decap_12
X_6068_ _6068_/A _6208_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_85_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_676 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1225 VGND VPWR sky130_fd_sc_hd__decap_8
X_5019_ _4971_/X _4972_/X _4962_/X _4973_/X _5019_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_26_410 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1197 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_56 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_605 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_402 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_11 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_44 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_811 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1074 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_367 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_518 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_99 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_837 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_510 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_297 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_531 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_971 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_1031 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_1053 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1102 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1097 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1124 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_825 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_911 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1146 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_313 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_741 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_711 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_593 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_755 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1062 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_668 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_145_359 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_679 VGND VPWR sky130_fd_sc_hd__decap_12
X_5370_ _4467_/A _4493_/X _5370_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_59_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_713 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_329 VGND VPWR sky130_fd_sc_hd__decap_6
X_4321_ _4310_/X _4314_/X _4310_/X _4314_/X _4321_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_4252_ _4252_/A _4253_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_7040_ _7040_/A _7040_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_113_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_407 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1191 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_4183_ _4847_/B _4459_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_68_844 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1172 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_941 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1055 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_387 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_847 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_1208 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_796 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_947 VGND VPWR sky130_fd_sc_hd__decap_6
X_6824_ _6822_/Y _6824_/B _6824_/X VGND VPWR sky130_fd_sc_hd__and2_4
XPHY_2209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_221 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_295 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_716 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_749 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1102 VGND VPWR sky130_fd_sc_hd__decap_6
X_6755_ _6744_/A _6744_/B _6744_/X _6754_/X _6804_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XPHY_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3967_ _3911_/Y _3965_/A _6034_/B _3967_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_91_1184 VGND VPWR sky130_fd_sc_hd__decap_12
X_5706_ _5689_/X _5692_/X _5707_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_17_1266 VGND VPWR sky130_fd_sc_hd__decap_8
X_6686_ _7689_/Q la_data_in[23] _6623_/X _6686_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_3898_ wbs_dat_i[1] _3882_/X _3899_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_192_922 VGND VPWR sky130_fd_sc_hd__decap_12
X_5637_ _5623_/X _5626_/X _5637_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_136_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_819 VGND VPWR sky130_fd_sc_hd__decap_4
X_5568_ _5325_/X _5326_/X _5298_/X _5327_/X _5568_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_151_318 VGND VPWR sky130_fd_sc_hd__decap_12
X_7307_ _3846_/X _7293_/X _7306_/X _7307_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_145_893 VGND VPWR sky130_fd_sc_hd__decap_12
X_4519_ _4519_/A _4485_/B _4519_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_176_1061 VGND VPWR sky130_fd_sc_hd__decap_6
X_5499_ _5464_/X _5478_/X _5464_/X _5478_/X _5499_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_160_841 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1045 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_554 VGND VPWR sky130_fd_sc_hd__decap_3
X_7238_ _7238_/A _7238_/B _7237_/Y _7238_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_120_727 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_68 VGND VPWR sky130_fd_sc_hd__decap_12
X_7169_ _7169_/A _7169_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_24_1215 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1234 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_674 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_398 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_495 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_1191 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_346 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_56 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_903 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_774 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_4145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_262 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_543 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_1084 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_593 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_243 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_468 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_930 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_799 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_98 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_440 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1246 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_169_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_490 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_663 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_635 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_487 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1153 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1036 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_874 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1039 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_516 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_741 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1271 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_733 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_886 VGND VPWR sky130_fd_sc_hd__decap_12
X_4870_ _4868_/X _4869_/X _4868_/X _4869_/X _4870_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_4690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1179 VGND VPWR sky130_fd_sc_hd__fill_1
X_3821_ _5602_/A _3798_/B _3821_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_33_788 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_991 VGND VPWR sky130_fd_sc_hd__fill_1
X_6540_ _6522_/Y _6523_/Y _6539_/X _6541_/B VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_158_440 VGND VPWR sky130_fd_sc_hd__decap_12
X_3752_ _7812_/Q _4614_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_119_816 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_580 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_304 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1050 VGND VPWR sky130_fd_sc_hd__decap_12
X_6471_ _6433_/X _6469_/X _6470_/Y _6471_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_185_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1130 VGND VPWR sky130_fd_sc_hd__decap_12
X_5422_ _4695_/A _4498_/B _5422_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_173_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_318 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_1231 VGND VPWR sky130_fd_sc_hd__decap_3
X_5353_ _5340_/X _5344_/X _5343_/X _5353_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_154_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_906 VGND VPWR sky130_fd_sc_hd__decap_12
X_4304_ _4303_/X _4304_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_173_1245 VGND VPWR sky130_fd_sc_hd__decap_12
X_5284_ _5229_/X _5273_/X _5229_/X _5273_/X _5284_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_102_738 VGND VPWR sky130_fd_sc_hd__decap_12
X_7023_ _7637_/Q la_data_in[67] _6961_/X _7023_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_4235_ _3728_/X _4235_/B _4236_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_114_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_4166_ _4158_/X _4165_/X _4158_/X _4165_/X _4166_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_210_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_696 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_184 VGND VPWR sky130_fd_sc_hd__decap_6
X_4097_ _4069_/X _4096_/X _4104_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_71_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_691 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_839 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_349 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_311 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6807_ _6754_/X _6806_/X _6785_/X _6807_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XPHY_2039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1227 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_788 VGND VPWR sky130_fd_sc_hd__decap_12
X_7787_ _7787_/D _7315_/A _7785_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4999_ _4997_/X _4998_/X _4997_/X _4998_/X _4999_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_24 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_366 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_440 VGND VPWR sky130_fd_sc_hd__decap_4
X_6738_ _6736_/Y _6737_/Y _6736_/Y _6737_/Y _6738_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1074 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_473 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_315 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1044 VGND VPWR sky130_fd_sc_hd__decap_6
X_6669_ _7695_/Q la_data_in[29] _6605_/X _6669_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_104_1066 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_977 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_668 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_1088 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_605 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_785 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_616 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_893 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_626 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_103 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_690 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_906 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_147 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_928 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_169 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1106 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_1042 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_505 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_825 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1113 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_696 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1139 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_633 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_292 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1179 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_733 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_300 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_26 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_788 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_276 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1130 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_736 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_760 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_922 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_972 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_281 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1098 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_936 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_318 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_969 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_852 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_405 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1017 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_909 VGND VPWR sky130_fd_sc_hd__decap_6
X_4020_ _4583_/A _4122_/B _4020_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_78_983 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_603 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_379 VGND VPWR sky130_fd_sc_hd__fill_1
X_5971_ _5967_/X _5968_/X _5974_/B _5972_/B VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_65_699 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_176 VGND VPWR sky130_fd_sc_hd__decap_8
X_7710_ _6567_/X _6498_/A _7707_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_198 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_593 VGND VPWR sky130_fd_sc_hd__decap_4
X_4922_ _4913_/X _4921_/X _4913_/X _4921_/X _4922_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_52_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1060 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_171 VGND VPWR sky130_fd_sc_hd__decap_12
X_7641_ _7015_/X _6947_/A _7624_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_205_1208 VGND VPWR sky130_fd_sc_hd__decap_12
X_4853_ _4016_/A _4854_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_33_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1077 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1230 VGND VPWR sky130_fd_sc_hd__decap_12
X_3804_ _5130_/A _4461_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_178_579 VGND VPWR sky130_fd_sc_hd__fill_1
X_7572_ _7572_/HI la_data_out[99] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_14_1203 VGND VPWR sky130_fd_sc_hd__decap_12
X_4784_ _4768_/X _4774_/X _4768_/X _4774_/X _4784_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1274 VGND VPWR sky130_fd_sc_hd__decap_3
X_6523_ la_data_in[4] _6523_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_146_410 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_1233 VGND VPWR sky130_fd_sc_hd__decap_12
X_3735_ _4829_/A _4479_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_20_279 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1258 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1217 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_679 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_27 VGND VPWR sky130_fd_sc_hd__decap_12
X_6454_ _7726_/Q la_data_in[124] _6390_/X _6454_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_162_914 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_498 VGND VPWR sky130_fd_sc_hd__fill_2
X_5405_ _5405_/A _5404_/X _5405_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_6385_ _7727_/Q _6387_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_133_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_703 VGND VPWR sky130_fd_sc_hd__decap_12
X_5336_ _5271_/X _5272_/X _5271_/X _5272_/X _5336_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_125_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_5267_ _5252_/X _5258_/X _5265_/X _5266_/X _5267_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_173_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_257 VGND VPWR sky130_fd_sc_hd__decap_12
X_7006_ _6982_/X _7005_/X _6999_/X _7006_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_102_568 VGND VPWR sky130_fd_sc_hd__decap_12
X_4218_ _4553_/A _4218_/B _4219_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_5198_ _5198_/A _3938_/A _5198_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_68_471 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_482 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_942 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_324 VGND VPWR sky130_fd_sc_hd__decap_12
X_4149_ _4111_/X _4141_/X _4142_/X _4148_/X _4149_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_28_346 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_143 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_474 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_609 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1194 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_23 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1002 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_552 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_703 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_855 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_747 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1008 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_11_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X _7746_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_911 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_398 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_966 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_165_763 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_445 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_20 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_479 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_769 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_460 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_666 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1082 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_658 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1274 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1116 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_179 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_3071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_371 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_141 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_686 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_387 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_944 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_730 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1105 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_903 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_454 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_762 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_711 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_6170_ _6167_/Y _6168_/X _6169_/X _7775_/D VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_170_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_682 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1245 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_5121_ _5098_/X _5104_/X _5092_/X _5105_/X _5121_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_170_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_706 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_877 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_257 VGND VPWR sky130_fd_sc_hd__decap_12
X_5052_ _5052_/A _4959_/B _5052_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_111_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_920 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1234 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_227 VGND VPWR sky130_fd_sc_hd__decap_12
X_4003_ _4925_/B _4123_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_37_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_441 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_666 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_923 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_485 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1008 VGND VPWR sky130_fd_sc_hd__decap_12
X_5954_ _5943_/X _5949_/X _5950_/X _5954_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_111_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_861 VGND VPWR sky130_fd_sc_hd__decap_12
X_4905_ _4902_/X _4903_/X _4904_/X _4905_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_40_319 VGND VPWR sky130_fd_sc_hd__decap_12
X_5885_ _5859_/X _5878_/B _5878_/X _5885_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_179_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1174 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_1005 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1185 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_522 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_708 VGND VPWR sky130_fd_sc_hd__decap_12
X_7624_ _7624_/D _7058_/A _7624_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_205_1038 VGND VPWR sky130_fd_sc_hd__decap_12
X_4836_ _4826_/X _4835_/X _4826_/X _4835_/X _4836_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_194_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1191 VGND VPWR sky130_fd_sc_hd__decap_12
X_7555_ _7555_/HI la_data_out[82] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_53_1082 VGND VPWR sky130_fd_sc_hd__decap_12
X_4767_ _4739_/X _4754_/X _4765_/X _4766_/X _4767_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_135_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1055 VGND VPWR sky130_fd_sc_hd__decap_12
X_6506_ _6504_/Y _6505_/Y _6506_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_193_379 VGND VPWR sky130_fd_sc_hd__decap_12
X_3718_ _3718_/A _4821_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_146_251 VGND VPWR sky130_fd_sc_hd__decap_12
X_7486_ _7486_/HI la_data_out[13] VGND VPWR sky130_fd_sc_hd__conb_1
X_4698_ _4698_/A _4698_/B _4698_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_107_638 VGND VPWR sky130_fd_sc_hd__decap_12
X_6437_ _6399_/X _6464_/B _6465_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_161_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1189 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_916 VGND VPWR sky130_fd_sc_hd__fill_1
X_6368_ _6354_/A _6368_/B _6368_/C _7734_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_0_404 VGND VPWR sky130_fd_sc_hd__decap_8
X_5319_ _4752_/X _4753_/X _4752_/X _4753_/X _5319_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_88_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_855 VGND VPWR sky130_fd_sc_hd__decap_12
X_6299_ _5975_/X _6299_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_130_674 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_611 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_931 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1059 VGND VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_2_1_1_wb_clk_i clkbuf_2_1_1_wb_clk_i/A clkbuf_3_3_0_wb_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_72_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_444 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_300 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_129 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_311 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_322 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_333 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_344 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_382 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_355 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_366 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_377 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_388 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_696 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_398 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_399 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1160 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_678 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_752 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_710 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_9 _6256_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_153_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_308 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_522 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_286 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_706 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_663 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_503 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_920 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_696 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_993 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_709 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1243 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_452 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_411 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_146 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_680 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_853 VGND VPWR sky130_fd_sc_hd__fill_1
X_5670_ _5668_/X _5669_/X _5668_/X _5669_/X _5670_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_176_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_864 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_1085 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_696 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1047 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_886 VGND VPWR sky130_fd_sc_hd__decap_12
X_4621_ _4603_/X _4620_/X _4603_/X _4620_/X _4621_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_124_1069 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_1060 VGND VPWR sky130_fd_sc_hd__decap_8
X_7340_ _7340_/A _7351_/B _7340_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_175_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_700 VGND VPWR sky130_fd_sc_hd__fill_2
X_4552_ _4552_/A _4595_/B _4552_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_204_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_593 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_744 VGND VPWR sky130_fd_sc_hd__decap_12
X_7271_ _7270_/Y _7265_/X _7271_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_171_530 VGND VPWR sky130_fd_sc_hd__decap_12
X_4483_ _5301_/B _4562_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_143_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_457 VGND VPWR sky130_fd_sc_hd__fill_1
X_6222_ _6219_/X _6220_/X _6221_/X _7766_/D VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_171_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_799 VGND VPWR sky130_fd_sc_hd__fill_1
X_6153_ _5050_/B _6152_/X _6020_/Y _6153_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_97_341 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_803 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1037 VGND VPWR sky130_fd_sc_hd__decap_12
X_5104_ _5099_/X _5103_/X _5102_/X _5104_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_44_1059 VGND VPWR sky130_fd_sc_hd__decap_8
X_6084_ _6158_/A _6084_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_112_685 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_525 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_216 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_184 VGND VPWR sky130_fd_sc_hd__decap_12
X_5035_ _4947_/X _4950_/Y _4952_/X _5035_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_100_869 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_27 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_4508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_928 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_3818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_978 VGND VPWR sky130_fd_sc_hd__decap_12
X_6986_ _6929_/Y _6931_/B _6931_/X _6985_/X _6986_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XPHY_3829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1111 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_5937_ _5931_/X _5934_/X _5935_/Y _5936_/X _5937_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_202_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1201 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_691 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_330 VGND VPWR sky130_fd_sc_hd__fill_2
X_5868_ _5865_/X _5866_/X _5865_/X _5866_/X _5868_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_210_943 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_864 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_341 VGND VPWR sky130_fd_sc_hd__decap_12
X_7607_ _7607_/D _7169_/A _7729_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_193_110 VGND VPWR sky130_fd_sc_hd__decap_12
X_4819_ _4630_/X _4636_/X _4623_/X _4637_/X _4819_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_210_976 VGND VPWR sky130_fd_sc_hd__decap_12
X_5799_ _5785_/X _5791_/X _5785_/X _5791_/X _5799_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_194_677 VGND VPWR sky130_fd_sc_hd__decap_12
X_7538_ _7538_/HI la_data_out[65] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_135_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_947 VGND VPWR sky130_fd_sc_hd__decap_12
X_7469_ _7469_/HI io_out[34] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_190_861 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_652 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_779 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1060 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_102 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_422 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_1025 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_764 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_130 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_803 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_141 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_611 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_163 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_824 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_174 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_185 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_312 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_196 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_683 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_346 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_356 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_379 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_711 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_733 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_850 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1023 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1026 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1250 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_799 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_939 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_812 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_385 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_845 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1051 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_923 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_422 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1095 VGND VPWR sky130_fd_sc_hd__decap_12
X_6840_ _6840_/A _6840_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_78_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_978 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1008 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_707 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_274 VGND VPWR sky130_fd_sc_hd__fill_1
X_6771_ _6709_/Y _6710_/Y _6770_/X _6771_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_165_1158 VGND VPWR sky130_fd_sc_hd__fill_1
X_3983_ _3971_/X _3982_/Y _3997_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_5722_ _5722_/A _5722_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_175_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_633 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_335 VGND VPWR sky130_fd_sc_hd__fill_1
X_5653_ _5651_/X _5652_/X _5651_/X _5652_/X _5653_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_4604_ _4820_/B _5300_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_176_688 VGND VPWR sky130_fd_sc_hd__decap_12
X_5584_ _5566_/X _5583_/X _5584_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_191_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1142 VGND VPWR sky130_fd_sc_hd__decap_12
X_7323_ io_in[16] _7323_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_11_1036 VGND VPWR sky130_fd_sc_hd__fill_1
X_4535_ _4535_/A _4793_/B _4535_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_132_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_27 VGND VPWR sky130_fd_sc_hd__decap_12
X_7254_ _7253_/X _7354_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_4466_ _4631_/B _4595_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_116_276 VGND VPWR sky130_fd_sc_hd__decap_12
X_6205_ _6189_/A _6205_/B _6205_/C _6207_/A VGND VPWR sky130_fd_sc_hd__nor3_4
X_7185_ _7245_/A _7184_/X _7246_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_4397_ _4392_/X _4396_/X _4395_/X _4397_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_131_257 VGND VPWR sky130_fd_sc_hd__decap_12
X_6136_ _4450_/X _6138_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_100_600 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_994 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_471 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_171 VGND VPWR sky130_fd_sc_hd__decap_12
X_6067_ _7327_/A _6063_/X _6066_/Y _6067_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_133_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_208 VGND VPWR sky130_fd_sc_hd__decap_12
X_5018_ _5000_/X _5001_/X _5000_/X _5001_/X _5018_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_100_688 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_794 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_293 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_4327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_989 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_3626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_466 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_617 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_414 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_769 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6969_ _7030_/A _6968_/X _6969_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_2925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_149 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_600 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_23 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_324 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_193 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1231 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_722 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_371 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_691 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_543 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_672 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_565 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_576 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_587 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1065 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_306 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_322 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_867 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_709 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_923 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_1158 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_325 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_967 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_791 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1074 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_672 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_992 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1044 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_636 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1107 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_891 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_861 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_703 VGND VPWR sky130_fd_sc_hd__decap_3
X_4320_ _4317_/X _4320_/B _6025_/C VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_154_894 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_425 VGND VPWR sky130_fd_sc_hd__fill_2
X_4251_ _4251_/A _4250_/X _4252_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_180_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_257 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1121 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_812 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_419 VGND VPWR sky130_fd_sc_hd__decap_8
X_4182_ _4182_/A _4847_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_79_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1067 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_517 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_851 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_550 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_723 VGND VPWR sky130_fd_sc_hd__decap_8
X_6823_ la_data_in[61] _6824_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_51_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_728 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1250 VGND VPWR sky130_fd_sc_hd__fill_1
X_6754_ _6747_/A _6747_/B _6747_/X _6753_/X _6754_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XPHY_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_609 VGND VPWR sky130_fd_sc_hd__fill_1
X_3966_ _7321_/A _3966_/B _6034_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_211_559 VGND VPWR sky130_fd_sc_hd__decap_12
X_5705_ _5670_/X _5671_/X _5670_/X _5671_/X _5705_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_143_1253 VGND VPWR sky130_fd_sc_hd__decap_12
X_6685_ _6668_/A _6685_/B _6684_/Y _7690_/D VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_137_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1196 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_480 VGND VPWR sky130_fd_sc_hd__decap_8
X_3897_ _5216_/A _3897_/B _3899_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_148_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_5636_ _5632_/Y _5635_/X _5632_/Y _5635_/X _5636_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_192_934 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_349 VGND VPWR sky130_fd_sc_hd__decap_12
X_5567_ _5558_/X _5559_/X _5558_/X _5559_/X _5567_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_105_703 VGND VPWR sky130_fd_sc_hd__decap_12
X_7306_ _7304_/Y _7324_/B _7306_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4518_ _4485_/A _4479_/B _4518_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_104_202 VGND VPWR sky130_fd_sc_hd__decap_12
X_5498_ _5494_/X _5497_/X _5494_/X _5497_/X _5498_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7237_ _7237_/A _7237_/B _7237_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_4449_ _4449_/A _4448_/X _6027_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_160_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1221 VGND VPWR sky130_fd_sc_hd__decap_12
X_7168_ _7166_/Y _7168_/B _7168_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_98_480 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_642 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1276 VGND VPWR sky130_fd_sc_hd__fill_1
X_6119_ _6119_/A _6118_/X _7783_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_59_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1246 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_964 VGND VPWR sky130_fd_sc_hd__decap_12
X_7099_ la_data_in[95] _7098_/B _7099_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_111_1219 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_837 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_720 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_196 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_742 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_358 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_509 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1011 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_701 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1025 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_797 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_274 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_391 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_419 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_110 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_945 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_675 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_338 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1080 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_123 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_989 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1061 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_499 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1165 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_330 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_1157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1048 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_753 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_717 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_391 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_542 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3820_ _4653_/A _5602_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_162_1139 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_288 VGND VPWR sky130_fd_sc_hd__decap_4
X_3751_ _3769_/A _3751_/B _3750_/Y _3751_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_158_452 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_828 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_451 VGND VPWR sky130_fd_sc_hd__decap_8
X_6470_ _6433_/X _6469_/X _6455_/X _6470_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_201_592 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1062 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_495 VGND VPWR sky130_fd_sc_hd__fill_1
X_5421_ _4716_/A _4505_/B _5421_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_145_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_5352_ _5347_/X _5351_/X _5350_/X _5352_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_86_1243 VGND VPWR sky130_fd_sc_hd__decap_8
X_4303_ _4301_/X _4302_/X _4303_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_114_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_918 VGND VPWR sky130_fd_sc_hd__decap_12
X_5283_ _5279_/X _5282_/X _5279_/X _5282_/X _5283_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_142_886 VGND VPWR sky130_fd_sc_hd__decap_12
X_7022_ _7012_/A _7022_/B _7022_/C _7022_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_87_428 VGND VPWR sky130_fd_sc_hd__decap_12
X_4234_ _3720_/A _4137_/X _4236_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_4_71 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_642 VGND VPWR sky130_fd_sc_hd__decap_12
X_4165_ _4163_/X _4164_/X _4162_/X _4165_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_110_750 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_506 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_623 VGND VPWR sky130_fd_sc_hd__decap_12
X_4096_ _4070_/Y _4095_/X _4094_/X _4096_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_209_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1017 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_818 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_27 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_233 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6806_ _6742_/A la_data_in[35] _6744_/X _6806_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_211_323 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_227 VGND VPWR sky130_fd_sc_hd__decap_12
X_4998_ _4430_/A _4429_/X _4430_/X _4998_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_7786_ _6094_/Y _7310_/A _7746_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_586 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_428 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_36 VGND VPWR sky130_fd_sc_hd__decap_8
X_3949_ _3728_/X _3949_/B _3951_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_6737_ la_data_in[37] _6737_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_183_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_485 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_1086 VGND VPWR sky130_fd_sc_hd__decap_12
X_6668_ _6668_/A _6661_/X _6667_/Y _6668_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_109_327 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_422 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_647 VGND VPWR sky130_fd_sc_hd__decap_6
X_5619_ _5618_/A _5617_/X _5618_/X _5619_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_180_904 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_764 VGND VPWR sky130_fd_sc_hd__decap_4
X_6599_ _6668_/A _6596_/A _6598_/X _6599_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_124_308 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_797 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_144_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1062 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1032 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_450 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_984 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1054 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1125 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_678 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_369 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_306 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_211 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_840 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_745 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_3242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_312 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_862 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_288 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_748 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_603 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1044 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_911 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_934 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_444 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_948 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_691 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_864 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_704 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_417 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_1029 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_660 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_428 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_671 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_601 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_995 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_358 VGND VPWR sky130_fd_sc_hd__decap_8
X_5970_ _5969_/X _5974_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_46_881 VGND VPWR sky130_fd_sc_hd__decap_4
X_4921_ _4914_/X _4920_/X _4914_/X _4920_/X _4921_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_391 VGND VPWR sky130_fd_sc_hd__decap_12
X_4852_ _4769_/A _4852_/B _4852_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7640_ _7640_/D _6950_/A _7624_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_178_536 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_586 VGND VPWR sky130_fd_sc_hd__decap_12
X_3803_ _4625_/A _5130_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_7571_ _7571_/HI la_data_out[98] VGND VPWR sky130_fd_sc_hd__conb_1
X_4783_ _4780_/X _4782_/X _4780_/X _4782_/X _4783_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_1089 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_1242 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1215 VGND VPWR sky130_fd_sc_hd__decap_12
X_6522_ _7702_/Q _6522_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_3734_ _7814_/Q _4829_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_159_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1245 VGND VPWR sky130_fd_sc_hd__decap_6
X_6453_ _6441_/X _6451_/X _6452_/Y _6453_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_174_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_989 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_926 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_477 VGND VPWR sky130_fd_sc_hd__fill_1
X_5404_ _5348_/A _4757_/B _5404_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_134_628 VGND VPWR sky130_fd_sc_hd__decap_12
X_6384_ _6382_/Y _6383_/Y _6382_/Y _6383_/Y _6449_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_162_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1002 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_1130 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_1013 VGND VPWR sky130_fd_sc_hd__decap_12
X_5335_ _5283_/X _5284_/X _5283_/X _5284_/X _5335_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_126_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1046 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1005 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_385 VGND VPWR sky130_fd_sc_hd__decap_12
X_5266_ _5252_/X _5258_/X _5252_/X _5258_/X _5266_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_141_171 VGND VPWR sky130_fd_sc_hd__decap_12
X_7005_ _7644_/Q la_data_in[74] _6940_/X _7005_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_4217_ _4505_/A _4217_/B _4219_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_87_269 VGND VPWR sky130_fd_sc_hd__decap_12
X_5197_ _5185_/X _5189_/X _5185_/X _5189_/X _5197_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_29_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_623 VGND VPWR sky130_fd_sc_hd__decap_12
X_4148_ _4132_/X _4179_/A _3918_/X _4235_/B _4148_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_68_494 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_678 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1151 VGND VPWR sky130_fd_sc_hd__decap_8
X_4079_ _4077_/X _4078_/X _4076_/X _4079_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_141_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_497 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_520 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_564 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_715 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1099 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_759 VGND VPWR sky130_fd_sc_hd__decap_4
X_7769_ _7769_/D _7769_/Q _7769_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_934 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_271 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_947 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_424 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_457 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_886 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1040 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_388 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_472 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_623 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1050 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1094 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_892 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_812 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_147 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_851 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_171 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1128 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_383 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_698 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_208 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_742 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_956 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_781 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_764 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_550 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_1128 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_774 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_723 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_801 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_981 VGND VPWR sky130_fd_sc_hd__fill_2
X_5120_ _5061_/X _5119_/X _5061_/X _5119_/X _5120_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_170_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1268 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_1227 VGND VPWR sky130_fd_sc_hd__decap_12
X_5051_ _4807_/X _4884_/X _4991_/X _5050_/X _5051_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_69_269 VGND VPWR sky130_fd_sc_hd__decap_12
X_4002_ _4455_/B _4925_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_66_932 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_453 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_935 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_380 VGND VPWR sky130_fd_sc_hd__decap_12
X_5953_ _5950_/X _5952_/X _5950_/X _5952_/X _5953_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_168_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_300 VGND VPWR sky130_fd_sc_hd__decap_12
X_4904_ _4902_/X _4903_/X _4904_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_34_873 VGND VPWR sky130_fd_sc_hd__decap_12
X_5884_ _5880_/X _5881_/X _5880_/X _5881_/X _5884_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_895 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1017 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1239 VGND VPWR sky130_fd_sc_hd__decap_12
X_7623_ _7128_/X _7623_/Q _7797_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_209_1197 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_534 VGND VPWR sky130_fd_sc_hd__decap_12
X_4835_ _4833_/X _4834_/X _4833_/X _4834_/X _4835_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_60_191 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_837 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_1050 VGND VPWR sky130_fd_sc_hd__decap_12
X_4766_ _4739_/X _4754_/X _4739_/X _4754_/X _4766_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7554_ _7554_/HI la_data_out[81] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_147_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_1020 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_1094 VGND VPWR sky130_fd_sc_hd__decap_4
X_3717_ _3733_/A _3717_/B _3716_/Y _7817_/D VGND VPWR sky130_fd_sc_hd__nor3_4
X_6505_ la_data_in[10] _6505_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_7485_ _7485_/HI la_data_out[12] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_101_1015 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1067 VGND VPWR sky130_fd_sc_hd__fill_1
X_4697_ _4697_/A _4657_/B _4698_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_146_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_6436_ _6400_/Y _6401_/Y _6468_/B _6464_/B VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_136_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_918 VGND VPWR sky130_fd_sc_hd__decap_12
X_6367_ wbs_dat_i[4] _6364_/B _6368_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_162_789 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_970 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_672 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_683 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_416 VGND VPWR sky130_fd_sc_hd__decap_12
X_5318_ _5314_/X _5317_/X _5314_/X _5317_/X _5318_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6298_ _6211_/A _6298_/B _6298_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_130_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_556 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_449 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_867 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_35 VGND VPWR sky130_fd_sc_hd__decap_12
X_5249_ _5245_/X _5248_/X _5245_/X _5248_/X _5249_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_69_770 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1005 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_902 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_913 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_166 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_23 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_188 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_56 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1109 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_147 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_301 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_312 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_489 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_323 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_322 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_334 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_821 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_345 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_692 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_356 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_394 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_367 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_208 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_378 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_44 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_389 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1251 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_701 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_959 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_722 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_745 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_907 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_298 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_718 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_1099 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1009 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_291 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_965 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_768 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_423 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_648 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_754 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_930 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_821 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_837 VGND VPWR sky130_fd_sc_hd__decap_12
X_4620_ _4611_/X _4619_/X _4611_/X _4619_/X _4620_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_163_1097 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1223 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_358 VGND VPWR sky130_fd_sc_hd__decap_8
X_4551_ _4546_/X _4550_/X _4549_/X _4551_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_184_881 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_263 VGND VPWR sky130_fd_sc_hd__decap_12
X_7270_ io_in[7] _7270_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4482_ _4482_/A _5301_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_144_756 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_542 VGND VPWR sky130_fd_sc_hd__decap_6
X_6221_ _5534_/Y _6216_/X _6194_/X _6221_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_48_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_277 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_428 VGND VPWR sky130_fd_sc_hd__decap_6
X_6152_ _4991_/X _6151_/X _6016_/Y _6152_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_135_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1163 VGND VPWR sky130_fd_sc_hd__decap_12
X_5103_ _5100_/X _5102_/B _5102_/X _5103_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_6083_ _6317_/C _6158_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_100_815 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_1049 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_1188 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_697 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_837 VGND VPWR sky130_fd_sc_hd__decap_12
X_5034_ _4974_/X _4975_/X _4953_/X _4976_/X _5034_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_111_196 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1098 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1110 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_3808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_743 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6985_ _6934_/A _6934_/B _6934_/X _6984_/X _6985_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_53_456 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_26 VGND VPWR sky130_fd_sc_hd__decap_8
X_5936_ _5931_/X _5934_/X _5931_/X _5934_/X _5936_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_179_631 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1131 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1213 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_141 VGND VPWR sky130_fd_sc_hd__decap_12
X_5867_ _5867_/A _5867_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_139_517 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_876 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_353 VGND VPWR sky130_fd_sc_hd__decap_12
X_7606_ _7238_/X _7606_/Q _7729_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4818_ _4617_/X _4618_/X _4611_/X _4619_/X _4818_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_5798_ _5795_/X _5796_/X _5805_/B _5798_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_210_988 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_550 VGND VPWR sky130_fd_sc_hd__decap_12
X_7537_ _7537_/HI la_data_out[64] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_181_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_689 VGND VPWR sky130_fd_sc_hd__decap_12
X_4749_ _4749_/A _4455_/B _4749_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_107_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_959 VGND VPWR sky130_fd_sc_hd__decap_12
X_7468_ _7468_/HI io_out[33] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_190_873 VGND VPWR sky130_fd_sc_hd__decap_12
X_6419_ la_data_in[114] _6420_/B VGND VPWR sky130_fd_sc_hd__inv_8
X_7399_ _7398_/Y _7387_/A _4434_/A _7257_/X wbs_dat_o[30] VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_150_737 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_202 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_973 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_984 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_472 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_686 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1010 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_740 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1072 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_710 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_637 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_114 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1015 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_787 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_106 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_120 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_142 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_815 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_153 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_164 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_814 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_175 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_836 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_186 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_695 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_818 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_870 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_368 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_572 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_391 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_1016 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_1035 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_618 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1038 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_552 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_428 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_394 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_375 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_209 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_1063 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_935 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_0 VGND VPWR sky130_fd_sc_hd__decap_3
X_3982_ _3914_/A _3999_/A _3981_/X _3979_/Y _3980_/Y _3982_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
X_6770_ _6770_/A _6769_/X _6770_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_35_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_106 VGND VPWR sky130_fd_sc_hd__decap_12
X_5721_ _5677_/X _5721_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_188_450 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_218 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_281 VGND VPWR sky130_fd_sc_hd__decap_12
X_5652_ _5503_/Y _5504_/X _5503_/Y _5504_/X _5652_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_206_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_684 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1151 VGND VPWR sky130_fd_sc_hd__decap_8
X_4603_ _4594_/X _4600_/X _4601_/X _4602_/X _4603_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_5583_ _5576_/X _5582_/X _5583_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_163_306 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_712 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_723 VGND VPWR sky130_fd_sc_hd__decap_8
X_4534_ _5294_/B _4793_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_7322_ _7370_/A _7322_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_144_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1211 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_907 VGND VPWR sky130_fd_sc_hd__decap_8
X_4465_ _4182_/A _4631_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_7253_ wbs_adr_i[2] _7253_/B _7253_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_172_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_715 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_726 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_288 VGND VPWR sky130_fd_sc_hd__decap_12
X_6204_ _5549_/X _6202_/Y _6205_/C VGND VPWR sky130_fd_sc_hd__nor2_4
X_7184_ _7181_/Y _7182_/Y _7181_/Y _7182_/Y _7184_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_113_940 VGND VPWR sky130_fd_sc_hd__decap_8
X_4396_ _4393_/X _4394_/X _4395_/X _4396_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_6135_ _6185_/A _6135_/B _7780_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_131_269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_973 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_835 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_623 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_27 VGND VPWR sky130_fd_sc_hd__decap_12
X_6066_ _7327_/A _6063_/X _7404_/A _6066_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_61_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_367 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_507 VGND VPWR sky130_fd_sc_hd__fill_1
X_5017_ _5006_/X _5007_/X _5006_/X _5007_/X _5017_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_261 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_434 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_4339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_562 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_629 VGND VPWR sky130_fd_sc_hd__decap_12
X_6968_ _6965_/Y _6966_/Y _6965_/Y _6966_/Y _6968_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_2915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_719 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_426 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5919_ _4742_/A _4532_/A _5919_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_2948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_107_1021 VGND VPWR sky130_fd_sc_hd__fill_1
X_6899_ _6875_/X _6897_/X _6898_/Y _7660_/D VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_146_1081 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1243 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_383 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_556 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_312 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_1077 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_838 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_721 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_592 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_242 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_779 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_741 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_420 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_644 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_648 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_198 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_873 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1081 VGND VPWR sky130_fd_sc_hd__fill_2
X_4250_ _4213_/X _4247_/X _4248_/Y _4249_/X _4250_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_45_1133 VGND VPWR sky130_fd_sc_hd__decap_12
X_4181_ _7737_/Q _4182_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_121_280 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_857 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_337 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_776 VGND VPWR sky130_fd_sc_hd__decap_12
X_6822_ _6822_/A _6822_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_23_426 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_757 VGND VPWR sky130_fd_sc_hd__decap_12
X_6753_ _6748_/Y _6749_/Y _6815_/B _6753_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_3965_ _3965_/A _3966_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_177_932 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_971 VGND VPWR sky130_fd_sc_hd__decap_12
X_5704_ _5679_/X _5704_/B _5704_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_104_1205 VGND VPWR sky130_fd_sc_hd__decap_12
X_3896_ _5341_/A _5216_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_6684_ _6620_/X _6684_/B _6684_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_143_1265 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_818 VGND VPWR sky130_fd_sc_hd__decap_12
X_5635_ _5633_/X _5634_/X _5633_/X _5634_/X _5635_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_148_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1249 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_391 VGND VPWR sky130_fd_sc_hd__decap_12
X_5566_ _5549_/X _5565_/X _5566_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_163_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1071 VGND VPWR sky130_fd_sc_hd__decap_12
X_7305_ _7276_/A _7324_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_4517_ _4512_/X _4516_/X _4515_/X _4517_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_160_810 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_489 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_715 VGND VPWR sky130_fd_sc_hd__decap_12
X_5497_ _5495_/X _5496_/X _5495_/X _5496_/X _5497_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_534 VGND VPWR sky130_fd_sc_hd__decap_12
X_7236_ _7238_/A _7236_/B _7236_/C _7607_/D VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_137_1036 VGND VPWR sky130_fd_sc_hd__fill_1
X_4448_ _6025_/C _4446_/Y _4318_/X _4447_/Y _4448_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_208_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_802 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1069 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_1233 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_898 VGND VPWR sky130_fd_sc_hd__decap_6
X_4379_ _4376_/Y _4378_/B _4378_/X _4379_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_7167_ la_data_in[102] _7168_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_150_1203 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_846 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_420 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_492 VGND VPWR sky130_fd_sc_hd__decap_8
X_6118_ _4038_/Y _6117_/X _6085_/X _6118_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_7098_ la_data_in[95] _7098_/B _7100_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_59_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_816 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_518 VGND VPWR sky130_fd_sc_hd__fill_1
X_6049_ _3910_/Y _6048_/X _6049_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_73_326 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_540 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_754 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_916 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1181 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1079 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1023 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_437 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_223 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_729 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_245 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1215 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_954 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_571 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1070 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_520 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_687 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_968 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_840 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1092 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1130 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_501 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_523 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_1125 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1177 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1008 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_353 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_624 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_337 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_18_732 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_1240 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_80 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_729 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_3980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_971 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3750_ wbs_dat_i[19] _3715_/X _3750_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_186_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_902 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_475 VGND VPWR sky130_fd_sc_hd__decap_12
X_5420_ _5420_/A _4497_/B _5420_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_199_1074 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_851 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_1154 VGND VPWR sky130_fd_sc_hd__decap_12
X_5351_ _5348_/X _5349_/X _5350_/X _5351_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_173_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_117 VGND VPWR sky130_fd_sc_hd__decap_12
X_4302_ _4283_/X _4284_/X _4282_/X _4285_/X _4302_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_126_394 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_691 VGND VPWR sky130_fd_sc_hd__decap_8
X_5282_ _5280_/X _5281_/X _5280_/X _5281_/X _5282_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_556 VGND VPWR sky130_fd_sc_hd__decap_12
X_4233_ _4215_/X _4232_/X _4215_/X _4232_/X _4233_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7021_ _7021_/A _7021_/B _7022_/C VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_142_898 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_83 VGND VPWR sky130_fd_sc_hd__decap_8
X_4164_ _4503_/A _4164_/B _4164_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_96_963 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_654 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_315 VGND VPWR sky130_fd_sc_hd__decap_12
X_4095_ _4092_/X _4093_/X _4094_/X _4095_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_56_849 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1029 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_540 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1004 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1207 VGND VPWR sky130_fd_sc_hd__decap_12
X_6805_ _6795_/A _6756_/X _6804_/Y _6805_/X VGND VPWR sky130_fd_sc_hd__and3_4
XPHY_2019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_919 VGND VPWR sky130_fd_sc_hd__decap_12
X_7785_ _7785_/D _7303_/A _7785_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4997_ _4964_/X _4965_/X _4963_/X _4966_/X _4997_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XPHY_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_335 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_239 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_56_1081 VGND VPWR sky130_fd_sc_hd__decap_12
X_6736_ _7671_/Q _6736_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_51_598 VGND VPWR sky130_fd_sc_hd__decap_12
X_3948_ _3935_/Y _3942_/X _3935_/Y _3942_/X _3948_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_139_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_6667_ _6602_/X _6667_/B _6667_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_139_59 VGND VPWR sky130_fd_sc_hd__fill_2
X_3879_ _5234_/A _5185_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_109_339 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_220 VGND VPWR sky130_fd_sc_hd__decap_12
X_5618_ _5618_/A _5617_/X _5618_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_6598_ _7698_/Q la_data_in[0] _6598_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_180_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_810 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1276 VGND VPWR sky130_fd_sc_hd__fill_1
X_5549_ _5547_/Y _5548_/X _5549_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_132_353 VGND VPWR sky130_fd_sc_hd__decap_12
X_7219_ _7199_/X _7218_/X _7212_/X _7219_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_154_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1074 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_56 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_996 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_304 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_529 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1066 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_318 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_562 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_342 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_814 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_690 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_532 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_324 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_548 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_740 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_32 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1143 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_32 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_615 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1029 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_996 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_851 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_990 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_372 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_832 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_459 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_342 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_6_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/A clkbuf_3_6_0_wb_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_97_716 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_749 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1261 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_1185 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1275 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1158 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_808 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_627 VGND VPWR sky130_fd_sc_hd__decap_12
X_4920_ _4918_/X _4919_/X _4918_/X _4919_/X _4920_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1013 VGND VPWR sky130_fd_sc_hd__decap_12
X_4851_ _4054_/A _4852_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_205_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_885 VGND VPWR sky130_fd_sc_hd__decap_8
X_3802_ _7806_/Q _4625_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_33_598 VGND VPWR sky130_fd_sc_hd__decap_12
X_7570_ _7570_/HI la_data_out[97] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_215 VGND VPWR sky130_fd_sc_hd__decap_4
X_4782_ _4568_/A _4782_/B _4782_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_53_1254 VGND VPWR sky130_fd_sc_hd__decap_12
X_6521_ _6519_/Y _6520_/Y _6519_/Y _6520_/Y _6521_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_3733_ _3733_/A _3731_/X _3732_/Y _3733_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_186_570 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_626 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_220 VGND VPWR sky130_fd_sc_hd__decap_12
X_6452_ _6441_/X _6451_/X _7404_/A _6452_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_174_776 VGND VPWR sky130_fd_sc_hd__decap_12
X_5403_ _5234_/A _4758_/B _5405_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_162_938 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_670 VGND VPWR sky130_fd_sc_hd__fill_1
X_6383_ la_data_in[126] _6383_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_5334_ _5332_/X _5334_/B _6228_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_47_1025 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_971 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_727 VGND VPWR sky130_fd_sc_hd__decap_12
X_5265_ _5262_/X _5264_/B _5274_/B _5265_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_134_1017 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_835 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_7004_ _6983_/X _7002_/X _7003_/Y _7004_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_173_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1203 VGND VPWR sky130_fd_sc_hd__fill_1
X_4216_ _4163_/X _4164_/X _4163_/X _4164_/X _4216_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_5196_ _5191_/X _5192_/X _5191_/X _5192_/X _5196_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_18_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_4147_ _4461_/B _4235_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_29_849 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_281 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_635 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_48 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_27 VGND VPWR sky130_fd_sc_hd__decap_12
X_4078_ _5294_/A _4078_/B _4078_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_43_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_532 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1045 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_312 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_576 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7768_ _6211_/Y _4540_/A _7769_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1179 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_507 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_187 VGND VPWR sky130_fd_sc_hd__decap_12
X_6719_ la_data_in[43] _6720_/B VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_570 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_208 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_760 VGND VPWR sky130_fd_sc_hd__decap_3
X_7699_ _6597_/X _6531_/A _7658_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_192_551 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_618 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_1040 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_489 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1204 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1136 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_469 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_602 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_484 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_944 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_925 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_871 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1221 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_532 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_86 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_154 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_395 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_557 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_581 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_220 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_754 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_968 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_253 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_1044 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_938 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_786 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1077 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_513 VGND VPWR sky130_fd_sc_hd__decap_12
X_5050_ _5050_/A _5050_/B _5050_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_170_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_1203 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_367 VGND VPWR sky130_fd_sc_hd__decap_12
X_4001_ _4641_/B _4455_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_78_771 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1113 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_808 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_465 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_605 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_156 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_95 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1264 VGND VPWR sky130_fd_sc_hd__decap_12
X_5952_ _5928_/X _5951_/X _5928_/X _5951_/X _5952_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_80_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_392 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_471 VGND VPWR sky130_fd_sc_hd__decap_12
X_4903_ _4479_/A _4903_/B _4903_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_5883_ _5858_/X _5988_/B _5883_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_178_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_502 VGND VPWR sky130_fd_sc_hd__decap_8
X_7622_ _7130_/X _7064_/A _7754_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4834_ _4612_/X _4616_/X _4615_/X _4834_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_179_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1029 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_546 VGND VPWR sky130_fd_sc_hd__decap_3
X_7553_ _7553_/HI la_data_out[80] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_159_570 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1062 VGND VPWR sky130_fd_sc_hd__decap_8
X_4765_ _4761_/X _4764_/X _4761_/X _4764_/X _4765_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6504_ _7708_/Q _6504_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_3716_ wbs_dat_i[23] _3715_/X _3716_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_105_1174 VGND VPWR sky130_fd_sc_hd__decap_12
X_7484_ _7484_/HI la_data_out[11] VGND VPWR sky130_fd_sc_hd__conb_1
X_4696_ _4680_/A _4666_/B _4698_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_135_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1253 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_1027 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1038 VGND VPWR sky130_fd_sc_hd__decap_12
X_6435_ _6467_/A _6467_/B _6468_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_175_1106 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_990 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_245 VGND VPWR sky130_fd_sc_hd__decap_12
X_6366_ _4366_/B _6373_/B _6368_/B VGND VPWR sky130_fd_sc_hd__and2_4
X_5317_ _5315_/X _5316_/X _5315_/X _5316_/X _5317_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_428 VGND VPWR sky130_fd_sc_hd__decap_6
X_6297_ _5980_/X _6073_/X _6296_/Y _5894_/A _6084_/X _6298_/B VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_130_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_568 VGND VPWR sky130_fd_sc_hd__decap_12
X_5248_ _5246_/X _5247_/X _5246_/X _5247_/X _5248_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_25_1120 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_47 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1191 VGND VPWR sky130_fd_sc_hd__decap_12
X_5179_ _5177_/X _5178_/X _5179_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_57_944 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_808 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_785 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_830 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_159 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_302 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_313 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_324 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_334 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_335 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_346 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_357 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_844 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_368 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_379 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_506 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_56 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1274 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_590 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_713 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_532 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_971 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_993 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1056 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_962 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_527 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_703 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_123 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_145 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_435 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_942 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1013 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_654 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_203_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1046 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_833 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_816 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_321 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_326 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_849 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1235 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_398 VGND VPWR sky130_fd_sc_hd__decap_6
X_4550_ _4549_/A _4549_/B _4549_/X _4550_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XPHY_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_916 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_927 VGND VPWR sky130_fd_sc_hd__decap_12
X_4481_ _4480_/Y _4482_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_6220_ _5582_/X _6199_/X _5582_/X _6199_/X _6220_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_143_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_407 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1142 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_289 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1093 VGND VPWR sky130_fd_sc_hd__decap_4
X_6151_ _6150_/X _6151_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_140_930 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1175 VGND VPWR sky130_fd_sc_hd__decap_12
X_5102_ _5100_/X _5102_/B _5102_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_6082_ _6189_/A _6080_/Y _6082_/C _6087_/A VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_83_1099 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_1069 VGND VPWR sky130_fd_sc_hd__decap_12
X_5033_ _5024_/X _5025_/X _5024_/X _5025_/X _5033_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_100_849 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_410 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_1055 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_711 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_722 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_733 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1050 VGND VPWR sky130_fd_sc_hd__decap_12
X_6984_ _6935_/Y _6937_/B _6937_/X _6983_/X _6984_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XPHY_3809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_755 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_137 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_780 VGND VPWR sky130_fd_sc_hd__decap_12
X_5935_ _7749_/Q _5935_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_80_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1143 VGND VPWR sky130_fd_sc_hd__decap_12
X_5866_ _5171_/A _4532_/A _5866_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_142_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_192 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1176 VGND VPWR sky130_fd_sc_hd__decap_12
X_7605_ _7241_/X _7605_/Q _7797_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4817_ _4810_/X _4816_/X _4810_/X _4816_/X _4817_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_107_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_365 VGND VPWR sky130_fd_sc_hd__fill_1
X_5797_ _5795_/X _5796_/X _5805_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_166_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_220 VGND VPWR sky130_fd_sc_hd__decap_12
X_7536_ _7536_/HI la_data_out[63] VGND VPWR sky130_fd_sc_hd__conb_1
X_4748_ _4455_/A _4748_/B _4748_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_147_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1050 VGND VPWR sky130_fd_sc_hd__decap_12
X_7467_ _7467_/HI io_out[32] VGND VPWR sky130_fd_sc_hd__conb_1
X_4679_ _4667_/A _4666_/B _4679_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_162_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_757 VGND VPWR sky130_fd_sc_hd__decap_12
X_6418_ _7716_/Q _6418_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_7398_ io_in[36] _7398_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_6349_ wbs_dat_i[9] _6349_/B _6349_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_88_310 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1215 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_855 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_996 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1022 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_752 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_722 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1084 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_126 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_799 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_44 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_110 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_118 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_121 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_440 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_143 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_321 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_602 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_855 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_154 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_945 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_422 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_176 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_849 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_187 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_326 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_674 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_198 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_848 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_668 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_551 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1071 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_882 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_245 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_705 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_779 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_1107 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1189 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_930 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_332 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_963 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1061 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1020 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_755 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1119 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1 VGND VPWR sky130_fd_sc_hd__decap_3
X_3981_ _3972_/X _3978_/X _3979_/Y _3980_/Y _3981_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_62_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_118 VGND VPWR sky130_fd_sc_hd__decap_12
X_5720_ _5678_/X _5717_/X _5718_/X _5719_/X _5722_/A VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_50_438 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_663 VGND VPWR sky130_fd_sc_hd__decap_8
X_5651_ _5647_/X _5648_/X _5649_/X _5650_/X _5651_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_203_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_123 VGND VPWR sky130_fd_sc_hd__decap_12
X_4602_ _4594_/X _4600_/X _4594_/X _4600_/X _4602_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_5582_ _5579_/A _5578_/X _5581_/Y _5582_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_141_1160 VGND VPWR sky130_fd_sc_hd__decap_12
X_7321_ _7321_/A _7321_/B _7321_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_163_329 VGND VPWR sky130_fd_sc_hd__decap_12
X_4533_ _5443_/B _5294_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_141_1193 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1253 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_532 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_94 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_391 VGND VPWR sky130_fd_sc_hd__decap_12
X_7252_ wbs_adr_i[1] wbs_adr_i[0] _7251_/Y _3709_/D _7253_/B VGND VPWR sky130_fd_sc_hd__or4_4
X_4464_ _4459_/X _4463_/X _4459_/X _4463_/X _4464_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6203_ _5549_/X _6202_/Y _6205_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_132_738 VGND VPWR sky130_fd_sc_hd__decap_6
X_7183_ _7602_/Q la_data_in[96] _7245_/A VGND VPWR sky130_fd_sc_hd__nand2_4
X_4395_ _4393_/X _4394_/X _4395_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_6134_ _6106_/X _6132_/X _6133_/X _7780_/Q _6109_/X _6135_/B VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_86_803 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_825 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_516 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_847 VGND VPWR sky130_fd_sc_hd__decap_12
X_6065_ _6068_/A _7404_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_133_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1150 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1101 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_1172 VGND VPWR sky130_fd_sc_hd__decap_12
X_5016_ _5005_/X _5009_/X _5005_/X _5009_/X _5016_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_27_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_755 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1219 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_777 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_917 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6967_ _6967_/A la_data_in[64] _7030_/A VGND VPWR sky130_fd_sc_hd__nand2_4
XPHY_3639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_585 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5918_ _5913_/X _5917_/X _5916_/X _5918_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XPHY_2938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_208 VGND VPWR sky130_fd_sc_hd__decap_12
X_6898_ _6875_/X _6897_/X _6811_/X _6898_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XPHY_2949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_635 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_972 VGND VPWR sky130_fd_sc_hd__decap_12
X_5849_ _5839_/X _5848_/X _5839_/X _5848_/X _5849_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_179_495 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_871 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_306 VGND VPWR sky130_fd_sc_hd__fill_2
X_7519_ _7519_/HI la_data_out[46] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_5_317 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_830 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_852 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_757 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_896 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_630 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_652 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1072 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1173 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1089 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_319 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1097 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_1048 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_733 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_424 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_703 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_574 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1111 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_1002 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_922 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1182 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1177 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_656 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_605 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_405 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_361 VGND VPWR sky130_fd_sc_hd__decap_12
X_4180_ _4179_/A _4179_/B _4179_/X _4180_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_122_760 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_1145 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_611 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_622 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_292 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_869 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_379 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_864 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_875 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_593 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_385 VGND VPWR sky130_fd_sc_hd__decap_12
X_6821_ _6819_/Y _6820_/Y _6819_/Y _6820_/Y _6821_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_169_1093 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_788 VGND VPWR sky130_fd_sc_hd__decap_8
X_6752_ _6814_/A _6814_/B _6815_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_3964_ _3963_/X _3965_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_211_528 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_769 VGND VPWR sky130_fd_sc_hd__decap_12
X_5703_ _5695_/X _5702_/X _5695_/X _5702_/X _5704_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_176_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_944 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1233 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_983 VGND VPWR sky130_fd_sc_hd__decap_12
X_6683_ _6668_/A _6655_/X _6682_/Y _6683_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_3895_ _5186_/A _5341_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_104_1217 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_977 VGND VPWR sky130_fd_sc_hd__decap_12
X_5634_ _4589_/A _5275_/X _5634_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_149_679 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_638 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_649 VGND VPWR sky130_fd_sc_hd__decap_12
X_5565_ _5550_/X _5564_/B _5564_/X _5565_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_157_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_532 VGND VPWR sky130_fd_sc_hd__decap_12
X_7304_ io_in[13] _7304_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_163_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1020 VGND VPWR sky130_fd_sc_hd__decap_3
X_4516_ _4515_/A _4514_/X _4515_/X _4516_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_89_1083 VGND VPWR sky130_fd_sc_hd__decap_12
X_5496_ _5432_/X _5433_/X _5432_/X _5433_/X _5496_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_145_885 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_502 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_727 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_7235_ _7235_/A _7190_/X _7236_/C VGND VPWR sky130_fd_sc_hd__nand2_4
X_4447_ _4447_/A _4447_/B _4447_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_132_546 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_719 VGND VPWR sky130_fd_sc_hd__decap_8
X_7166_ _7608_/Q _7166_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4378_ _4376_/Y _4378_/B _4378_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_86_622 VGND VPWR sky130_fd_sc_hd__decap_12
X_6117_ _6158_/A _6117_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_85_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_335 VGND VPWR sky130_fd_sc_hd__fill_1
X_7097_ io_out[5] _7096_/X _7098_/B VGND VPWR sky130_fd_sc_hd__xnor2_4
X_6048_ _6042_/A _3909_/Y _6058_/B _6048_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_160_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_891 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_338 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1025 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1160 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_861 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1005 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_552 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_766 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1069 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_703 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_928 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1193 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_8_0_wb_clk_i clkbuf_4_9_0_wb_clk_i/A _7729_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_3436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1035 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1068 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_235 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1199 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_922 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_257 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_281 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_752 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_633 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_318 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_699 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_852 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1096 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_1164 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_821 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_1137 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1189 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_320 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_365 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_688 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_880 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_636 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_206_812 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_850 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_202 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_747 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_410 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_933 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_983 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_914 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_487 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_159 VGND VPWR sky130_fd_sc_hd__decap_12
X_5350_ _5348_/X _5349_/X _5350_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_142_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1223 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_980 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1207 VGND VPWR sky130_fd_sc_hd__decap_12
X_4301_ _4301_/A _4301_/B _4301_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_160_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_5281_ _5059_/Y _5060_/X _5059_/Y _5060_/X _5281_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_257 VGND VPWR sky130_fd_sc_hd__decap_12
X_7020_ _7012_/A _6975_/X _7019_/Y _7020_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_141_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_568 VGND VPWR sky130_fd_sc_hd__decap_12
X_4232_ _4216_/X _4222_/X _4223_/X _4231_/X _4232_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_68_633 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_110 VGND VPWR sky130_fd_sc_hd__decap_12
X_4163_ _4162_/A _4161_/X _4162_/X _4163_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_136_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_953 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_975 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_452 VGND VPWR sky130_fd_sc_hd__decap_12
X_4094_ _4092_/X _4093_/X _4094_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_55_327 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_552 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_872 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_708 VGND VPWR sky130_fd_sc_hd__decap_12
X_6804_ _6741_/X _6804_/B _6804_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XPHY_2009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7784_ _7784_/D _7784_/Q _7746_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_180_1219 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_190 VGND VPWR sky130_fd_sc_hd__decap_12
X_4996_ _4956_/X _4957_/X _4958_/X _4959_/X _4996_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_23_257 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_408 VGND VPWR sky130_fd_sc_hd__decap_12
X_6735_ _6735_/A _6735_/B _6735_/X VGND VPWR sky130_fd_sc_hd__and2_4
XPHY_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3947_ _3943_/X _3946_/Y _3947_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_56_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1003 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_605 VGND VPWR sky130_fd_sc_hd__decap_4
X_6666_ _6885_/A _6666_/B _6665_/X _6666_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_176_251 VGND VPWR sky130_fd_sc_hd__decap_12
X_3878_ _4743_/A _5234_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_30_1200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1099 VGND VPWR sky130_fd_sc_hd__decap_12
X_5617_ _4718_/A _4613_/B _5617_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_104_1058 VGND VPWR sky130_fd_sc_hd__decap_8
X_6597_ _6668_/A _6535_/X _6597_/C _6597_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_191_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_928 VGND VPWR sky130_fd_sc_hd__decap_12
X_5548_ _5548_/A _5546_/X _5548_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_155_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_822 VGND VPWR sky130_fd_sc_hd__decap_12
X_5479_ _5420_/X _5424_/X _5420_/X _5424_/X _5479_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_155_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_855 VGND VPWR sky130_fd_sc_hd__decap_12
X_7218_ _7151_/A la_data_in[107] _7153_/X _7218_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_59_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_398 VGND VPWR sky130_fd_sc_hd__decap_12
X_7149_ la_data_in[108] _7150_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_113_590 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_785 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_316 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1078 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_349 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_56 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_574 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_354 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_544 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_886 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_752 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_44 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1155 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_881 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_44 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_928 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_427 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_384 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_630 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_877 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_728 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_931 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1273 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_452 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_1197 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_923 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_338 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_842 VGND VPWR sky130_fd_sc_hd__decap_12
X_4850_ _4839_/X _4849_/X _4839_/X _4849_/X _4850_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_72_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1025 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_196 VGND VPWR sky130_fd_sc_hd__decap_12
X_3801_ _3791_/A _3798_/X _3800_/Y _3801_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_159_730 VGND VPWR sky130_fd_sc_hd__fill_2
X_4781_ _4565_/B _4782_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_60_396 VGND VPWR sky130_fd_sc_hd__fill_1
X_6520_ la_data_in[5] _6520_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_140_1203 VGND VPWR sky130_fd_sc_hd__fill_2
X_3732_ wbs_dat_i[21] _3715_/X _3732_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_158_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_892 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_261 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_391 VGND VPWR sky130_fd_sc_hd__decap_12
X_6451_ _7727_/Q la_data_in[125] _6387_/X _6451_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_173_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_608 VGND VPWR sky130_fd_sc_hd__decap_12
X_5402_ _5072_/A _4756_/B _5402_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_174_788 VGND VPWR sky130_fd_sc_hd__decap_12
X_6382_ _7728_/Q _6382_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_5333_ _5332_/A _5331_/X _5334_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_115_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_983 VGND VPWR sky130_fd_sc_hd__decap_12
X_5264_ _5262_/X _5264_/B _5274_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_130_825 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_739 VGND VPWR sky130_fd_sc_hd__decap_12
X_7003_ _6983_/X _7002_/X _6999_/X _7003_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_141_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1029 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_398 VGND VPWR sky130_fd_sc_hd__decap_12
X_4215_ _4166_/X _4175_/X _4166_/X _4175_/X _4215_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_5195_ _5168_/X _5194_/X _5168_/X _5194_/X _5195_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_205_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_62 VGND VPWR sky130_fd_sc_hd__decap_12
X_4146_ _4758_/B _4461_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_60_1248 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_593 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_967 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_135 VGND VPWR sky130_fd_sc_hd__decap_8
X_4077_ _4074_/X _4075_/X _4076_/X _4077_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_141_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1035 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_341 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_886 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4979_ _4977_/X _4978_/X _4977_/X _4978_/X _4979_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7767_ _6218_/Y _7767_/Q _7769_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_829 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6718_ _6718_/A _6720_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_7698_ _6599_/X _7698_/Q _7658_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_211_199 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_733 VGND VPWR sky130_fd_sc_hd__decap_4
X_6649_ _6695_/A _6695_/B _6696_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_20_783 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_563 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_905 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1052 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_427 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_630 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_332 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1265 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1216 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_56 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_901 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_923 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_956 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_989 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_937 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_883 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_500 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_959 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_3030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_203_623 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1266 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_645 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_184 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_98 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_166 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_379 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_914 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_571 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_936 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_777 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_297 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_769 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_961 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1081 VGND VPWR sky130_fd_sc_hd__decap_3
X_4000_ _4000_/A _4641_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_111_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_783 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_135 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_1125 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_477 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_168 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_263 VGND VPWR sky130_fd_sc_hd__decap_12
X_5951_ _5938_/X _5940_/X _5951_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_52_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1276 VGND VPWR sky130_fd_sc_hd__fill_1
X_4902_ _4902_/A _5129_/B _4902_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_33_330 VGND VPWR sky130_fd_sc_hd__decap_12
X_5882_ _5878_/X _5879_/X _5880_/X _5881_/X _5988_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_206_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_672 VGND VPWR sky130_fd_sc_hd__decap_12
X_4833_ _4828_/X _4832_/X _4828_/X _4832_/X _4833_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7621_ _7133_/X _7621_/Q _7624_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_7552_ _7552_/HI la_data_out[79] VGND VPWR sky130_fd_sc_hd__conb_1
X_4764_ _4762_/X _4763_/X _4762_/X _4763_/X _4764_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_119_402 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1120 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_582 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1025 VGND VPWR sky130_fd_sc_hd__decap_8
X_6503_ _6503_/A _6502_/Y _6503_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_147_733 VGND VPWR sky130_fd_sc_hd__decap_4
X_3715_ _3759_/A _3715_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_147_744 VGND VPWR sky130_fd_sc_hd__decap_12
X_7483_ _7483_/HI la_data_out[10] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_179_1221 VGND VPWR sky130_fd_sc_hd__decap_12
X_4695_ _4695_/A _4665_/B _4695_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_105_1186 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_703 VGND VPWR sky130_fd_sc_hd__decap_12
X_6434_ _6403_/Y _6405_/B _6405_/X _6433_/X _6467_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_135_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1265 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_6365_ _6354_/A _6365_/B _6364_/Y _7735_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_161_257 VGND VPWR sky130_fd_sc_hd__decap_12
X_5316_ _5169_/X _5173_/X _5172_/X _5316_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_130_600 VGND VPWR sky130_fd_sc_hd__decap_12
X_6296_ _5953_/X _5979_/X _6296_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_103_836 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_15 VGND VPWR sky130_fd_sc_hd__fill_1
X_5247_ _5084_/X _5088_/X _5084_/X _5088_/X _5247_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_76_709 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_666 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_368 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1132 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_699 VGND VPWR sky130_fd_sc_hd__decap_3
X_5178_ _5178_/A _4743_/B _5178_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_111_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1067 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_956 VGND VPWR sky130_fd_sc_hd__decap_12
X_4129_ _4113_/X _4120_/X _4121_/X _4128_/X _4129_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_186_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1146 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_390 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_989 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_959 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_127 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_600 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_611 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_303 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_314 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_325 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_336 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_347 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_346 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_171 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_358 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_369 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_35 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_558 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_529 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_725 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_245 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_983 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_514 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_536 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_644 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1210 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_974 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_539 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_157 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_712 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_820 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_447 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_789 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_970 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_672 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_886 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_187_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_845 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_333 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1203 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_891 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_338 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_733 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1247 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_939 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_562 VGND VPWR sky130_fd_sc_hd__fill_2
X_4480_ _4480_/A _4480_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_128_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1091 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_257 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1121 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_419 VGND VPWR sky130_fd_sc_hd__decap_8
X_6150_ _4884_/X _6150_/B _6150_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_174_1162 VGND VPWR sky130_fd_sc_hd__decap_12
X_5101_ _5095_/A _5129_/B _5102_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_170_1015 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_333 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1187 VGND VPWR sky130_fd_sc_hd__decap_3
X_6081_ _6081_/A _6079_/X _6082_/C VGND VPWR sky130_fd_sc_hd__and2_4
Xclkbuf_4_10_0_wb_clk_i clkbuf_3_5_0_wb_clk_i/X _7785_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_57_208 VGND VPWR sky130_fd_sc_hd__decap_8
X_5032_ _5032_/A _5032_/B _5050_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_211_1067 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_550 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_764 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_561 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_403 VGND VPWR sky130_fd_sc_hd__decap_12
X_6983_ _6940_/A _6940_/B _6940_/X _6982_/X _6983_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_20_1062 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_149 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_767 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_190 VGND VPWR sky130_fd_sc_hd__decap_12
X_5934_ _5932_/X _5933_/X _5934_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_179_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1005 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_812 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_288 VGND VPWR sky130_fd_sc_hd__decap_12
X_5865_ _5863_/X _5864_/X _5862_/X _5865_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_167_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_480 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_1155 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_828 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1117 VGND VPWR sky130_fd_sc_hd__decap_12
X_4816_ _4811_/X _4815_/X _4811_/X _4815_/X _4816_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7604_ _7244_/X _7604_/Q _7729_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_166_316 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1188 VGND VPWR sky130_fd_sc_hd__decap_3
X_5796_ _4680_/A _4491_/A _5796_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_166_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_135 VGND VPWR sky130_fd_sc_hd__decap_12
X_4747_ _4747_/A _4747_/B _4747_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7535_ _7535_/HI la_data_out[62] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_119_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_27 VGND VPWR sky130_fd_sc_hd__decap_12
X_7466_ _7466_/HI io_out[31] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_134_202 VGND VPWR sky130_fd_sc_hd__decap_12
X_4678_ _4678_/A _4665_/B _4678_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_179_1062 VGND VPWR sky130_fd_sc_hd__decap_12
X_6417_ _6415_/Y _6417_/B _6417_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_162_544 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_769 VGND VPWR sky130_fd_sc_hd__decap_12
X_7397_ _7396_/Y _7387_/X _7775_/Q _7388_/X wbs_dat_o[29] VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6348_ _4235_/B _6348_/B _6350_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_88_300 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_322 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_953 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_644 VGND VPWR sky130_fd_sc_hd__decap_8
X_6279_ _5858_/X _5988_/B _5988_/X _6279_/Y VGND VPWR sky130_fd_sc_hd__a21boi_4
XFILLER_163_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_208 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1192 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1034 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_509 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_68 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_1044 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1096 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_447 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_138 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_239 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_100 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_672 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_122 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_56 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_133 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_480 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_452 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_155 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_333 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_867 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_177 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_636 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_957 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_434 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_188 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_1050 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_703 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1083 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_71 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1242 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_717 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_374 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_482 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_942 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_344 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_975 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_782 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_793 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1073 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_556 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_567 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_520 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_531 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_745 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_767 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_609 VGND VPWR sky130_fd_sc_hd__fill_1
X_3980_ _3978_/X _3980_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_2 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_806 VGND VPWR sky130_fd_sc_hd__decap_12
X_5650_ _5647_/X _5648_/X _5647_/X _5648_/X _5650_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_188_485 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_152 VGND VPWR sky130_fd_sc_hd__fill_1
X_4601_ _4552_/X _4556_/X _4555_/X _4601_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_148_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_135 VGND VPWR sky130_fd_sc_hd__decap_12
X_5581_ _5581_/A _5581_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_54_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_563 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1221 VGND VPWR sky130_fd_sc_hd__decap_12
X_7320_ _7259_/A _7321_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_141_1172 VGND VPWR sky130_fd_sc_hd__decap_4
X_4532_ _4532_/A _5443_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_190_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_820 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1265 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_0_1_wb_clk_i clkbuf_2_0_1_wb_clk_i/A clkbuf_2_0_1_wb_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_7251_ wbs_adr_i[3] _7251_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_171_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1178 VGND VPWR sky130_fd_sc_hd__decap_12
X_4463_ _4462_/A _4462_/B _4462_/X _4463_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_117_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1208 VGND VPWR sky130_fd_sc_hd__decap_12
X_6202_ _5564_/X _6202_/B _6202_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_7182_ la_data_in[97] _7182_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_113_920 VGND VPWR sky130_fd_sc_hd__fill_1
X_4394_ _4590_/A _4394_/B _4394_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_98_642 VGND VPWR sky130_fd_sc_hd__decap_12
X_6133_ _6123_/Y _6133_/B _6133_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_112_430 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_815 VGND VPWR sky130_fd_sc_hd__decap_8
X_6064_ wb_rst_i _6068_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_859 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_347 VGND VPWR sky130_fd_sc_hd__decap_12
X_5015_ _5012_/A _5013_/A _5014_/X _5032_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_61_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1203 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1225 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_285 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_391 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_3607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1217 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6966_ la_data_in[65] _6966_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_198_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_929 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_119 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_597 VGND VPWR sky130_fd_sc_hd__decap_12
X_5917_ _5914_/X _5915_/X _5916_/X _5917_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XPHY_2928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_452 VGND VPWR sky130_fd_sc_hd__decap_12
X_6897_ _7660_/Q la_data_in[58] _6833_/X _6897_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_210_721 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_642 VGND VPWR sky130_fd_sc_hd__decap_12
X_5848_ _5807_/Y _5808_/X _5807_/Y _5808_/X _5848_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_194_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_984 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_195_989 VGND VPWR sky130_fd_sc_hd__decap_12
X_5779_ _5776_/X _5777_/X _5778_/X _5779_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_182_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_883 VGND VPWR sky130_fd_sc_hd__fill_2
X_7518_ _7518_/HI la_data_out[45] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_5_329 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_190 VGND VPWR sky130_fd_sc_hd__decap_12
X_7449_ _7449_/HI io_out[14] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_190_650 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1130 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_642 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_664 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1084 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1095 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_1005 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_686 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1185 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_496 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_807 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1128 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_959 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1000 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_981 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_288 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1150 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_772 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_614 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_934 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1156 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_658 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1099 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_668 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_371 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_555 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1099 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_886 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_417 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_728 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_590 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_818 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_561 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_887 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_898 VGND VPWR sky130_fd_sc_hd__decap_12
X_6820_ la_data_in[62] _6820_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_24_929 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_575 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_277 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1111 VGND VPWR sky130_fd_sc_hd__decap_12
X_3963_ _3993_/A _3962_/X _3963_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_6751_ _6748_/Y _6749_/Y _6748_/Y _6749_/Y _6814_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_195_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1264 VGND VPWR sky130_fd_sc_hd__decap_12
X_5702_ _5700_/X _5701_/X _5700_/X _5701_/X _5702_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
Xclkbuf_1_1_0_wb_clk_i clkbuf_0_wb_clk_i/X clkbuf_1_1_0_wb_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_6682_ _6617_/X _6654_/X _6682_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_189_794 VGND VPWR sky130_fd_sc_hd__decap_12
X_3894_ _5787_/A _5186_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_176_422 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_956 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_995 VGND VPWR sky130_fd_sc_hd__decap_12
X_5633_ _5633_/A _5603_/X _5633_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_104_1229 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_989 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_191_403 VGND VPWR sky130_fd_sc_hd__decap_12
X_5564_ _5550_/X _5564_/B _5564_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_192_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_690 VGND VPWR sky130_fd_sc_hd__decap_12
X_4515_ _4515_/A _4514_/X _4515_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7303_ _7303_/A _7292_/B _7303_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_156_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_330 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_544 VGND VPWR sky130_fd_sc_hd__decap_4
X_5495_ _5474_/X _5475_/X _5471_/X _5476_/X _5495_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_89_1095 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_588 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_514 VGND VPWR sky130_fd_sc_hd__decap_4
X_4446_ _4385_/X _4444_/Y _4445_/X _4446_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
X_7234_ _6052_/A _7238_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_171_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_856 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1098 VGND VPWR sky130_fd_sc_hd__fill_2
X_7165_ _7163_/Y _7165_/B _7165_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_4377_ _4369_/X _4370_/X _4372_/X _4378_/B VGND VPWR sky130_fd_sc_hd__o21a_4
X_6116_ _6189_/A _6114_/Y _6116_/C _6119_/A VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_113_794 VGND VPWR sky130_fd_sc_hd__decap_6
X_7096_ _7034_/Y _7035_/Y _7095_/X _7096_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_86_634 VGND VPWR sky130_fd_sc_hd__decap_6
X_6047_ _6333_/A _6332_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_39_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_306 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_27 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_4105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_113_1082 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_520 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_1037 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_4116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_514 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_1044 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_873 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1017 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_406 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_709 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1178 VGND VPWR sky130_fd_sc_hd__decap_12
X_6949_ _6947_/Y _6949_/B _6949_/X VGND VPWR sky130_fd_sc_hd__and2_4
XPHY_2725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_951 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_400 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_269 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_511 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_148 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_661 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_672 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1274 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_1176 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1149 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_750 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_772 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_591 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_818 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_712 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_380 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1087 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_233 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_586 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_93 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_208 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_567 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_483 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_926 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1194 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_812 VGND VPWR sky130_fd_sc_hd__decap_12
X_4300_ _4824_/A _4299_/X _4301_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_173_1205 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_992 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_374 VGND VPWR sky130_fd_sc_hd__decap_12
X_5280_ _5268_/X _5269_/X _5267_/X _5270_/X _5280_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_153_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1219 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_30 VGND VPWR sky130_fd_sc_hd__fill_1
X_4231_ _4227_/X _4229_/X _4240_/B _4231_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_99_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_910 VGND VPWR sky130_fd_sc_hd__decap_12
X_4162_ _4162_/A _4161_/X _4162_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_136_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_764 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_987 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_464 VGND VPWR sky130_fd_sc_hd__decap_12
X_4093_ _4039_/X _4064_/X _4065_/X _4093_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_55_339 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_520 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_391 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_737 VGND VPWR sky130_fd_sc_hd__decap_12
X_6803_ _6795_/A _6758_/X _6802_/Y _7671_/D VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_211_304 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1081 VGND VPWR sky130_fd_sc_hd__decap_12
X_7783_ _7783_/D _7783_/Q _7746_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4995_ _4968_/X _4969_/X _4967_/X _4970_/X _4995_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_17_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_269 VGND VPWR sky130_fd_sc_hd__decap_12
X_6734_ la_data_in[38] _6735_/B VGND VPWR sky130_fd_sc_hd__inv_8
X_3946_ _3946_/A _3946_/B _3946_/Y VGND VPWR sky130_fd_sc_hd__xnor2_4
XFILLER_20_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_444 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_764 VGND VPWR sky130_fd_sc_hd__decap_12
X_3877_ _3877_/A _4743_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_6665_ la_data_in[31] _6663_/Y _6665_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_139_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_954 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1105 VGND VPWR sky130_fd_sc_hd__decap_12
X_5616_ _4743_/A _4291_/A _5618_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_30_1212 VGND VPWR sky130_fd_sc_hd__decap_12
X_6596_ _6596_/A _6596_/B _6597_/C VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_145_650 VGND VPWR sky130_fd_sc_hd__decap_12
X_5547_ _5548_/A _5546_/X _5547_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_145_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_620 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_834 VGND VPWR sky130_fd_sc_hd__decap_12
X_5478_ _5465_/X _5477_/X _5478_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_160_631 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_867 VGND VPWR sky130_fd_sc_hd__decap_12
X_4429_ _4426_/X _4428_/X _4425_/X _4429_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_7217_ _7200_/X _7215_/X _7216_/Y _7217_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_105_569 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1130 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_720 VGND VPWR sky130_fd_sc_hd__decap_12
X_7148_ _7614_/Q _7150_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_171_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1002 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_111 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1212 VGND VPWR sky130_fd_sc_hd__decap_8
X_7079_ _7070_/Y _7071_/Y _7072_/X _7078_/X _7079_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_171_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_328 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_147 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_810 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_586 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_154_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_208 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1150 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1120 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_589 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_781 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_56 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_893 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_291 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_712 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_936 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_959 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_864 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_341 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_439 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_685 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_943 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_807 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_935 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_692 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_597 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_707 VGND VPWR sky130_fd_sc_hd__decap_12
X_3800_ wbs_dat_i[13] _3822_/B _3800_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_4780_ _4779_/A _4779_/B _4779_/X _4780_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_207_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_206 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3731_ _4793_/A _3712_/X _3731_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_174_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_6450_ _6057_/A _6450_/B _6450_/C _7728_/D VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_147_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_273 VGND VPWR sky130_fd_sc_hd__decap_12
X_5401_ _5356_/X _5357_/X _5356_/X _5357_/X _5401_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6381_ _6381_/A _6381_/B _6381_/C _6381_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_103_1070 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1021 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_428 VGND VPWR sky130_fd_sc_hd__decap_12
X_5332_ _5332_/A _5331_/X _5332_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_114_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1038 VGND VPWR sky130_fd_sc_hd__decap_8
X_5263_ _4459_/A _4782_/B _5264_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_170_995 VGND VPWR sky130_fd_sc_hd__decap_12
X_4214_ _4177_/X _4192_/X _4177_/X _4192_/X _4214_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7002_ _7645_/Q la_data_in[75] _6937_/X _7002_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_5194_ _5183_/X _5193_/X _5183_/X _5193_/X _5194_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_141_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_431 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_1216 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_442 VGND VPWR sky130_fd_sc_hd__decap_12
X_4145_ _4145_/A _4758_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_56_615 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_74 VGND VPWR sky130_fd_sc_hd__decap_12
X_4076_ _4074_/X _4075_/X _4076_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_84_979 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_481 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1150 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_489 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_843 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_353 VGND VPWR sky130_fd_sc_hd__decap_12
X_7766_ _7766_/D _5534_/A _7769_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_898 VGND VPWR sky130_fd_sc_hd__decap_12
X_4978_ _4938_/X _4939_/X _4892_/X _4940_/X _4978_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XPHY_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_156 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6717_ _6717_/A _6717_/B _6717_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_177_550 VGND VPWR sky130_fd_sc_hd__decap_12
X_3929_ _4654_/A _3930_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_7697_ _6666_/Y io_out[1] _7696_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_138_926 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_520 VGND VPWR sky130_fd_sc_hd__decap_12
X_6648_ _6630_/Y _6631_/Y _6698_/B _6695_/B VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_166_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_795 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1020 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_575 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_917 VGND VPWR sky130_fd_sc_hd__decap_12
X_6579_ _7705_/Q la_data_in[7] _6515_/X _6579_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_106_812 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1064 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_981 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_416 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_439 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1105 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_951 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_344 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_729 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_751 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_919 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_114 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_294 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_968 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_602 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_62 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1207 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1215 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_3053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1237 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_657 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_196 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_178 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_881 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_93 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_892 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_733 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_918 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_789 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_575 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_70 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_973 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_815 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_314 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1041 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_795 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_851 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_93_776 VGND VPWR sky130_fd_sc_hd__decap_12
X_5950_ _5943_/X _5949_/X _5950_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_207_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_821 VGND VPWR sky130_fd_sc_hd__decap_3
X_4901_ _4901_/A _5129_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_80_459 VGND VPWR sky130_fd_sc_hd__decap_12
X_5881_ _5878_/X _5879_/X _5878_/X _5879_/X _5881_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_206_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_342 VGND VPWR sky130_fd_sc_hd__decap_12
X_7620_ _7620_/D _7070_/A _7624_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4832_ _4829_/X _4830_/X _4831_/X _4832_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_61_684 VGND VPWR sky130_fd_sc_hd__decap_12
X_7551_ _7551_/HI la_data_out[78] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_159_550 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_306 VGND VPWR sky130_fd_sc_hd__decap_12
X_4763_ _4467_/X _4471_/X _4467_/X _4471_/X _4763_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_119_414 VGND VPWR sky130_fd_sc_hd__decap_12
X_6502_ la_data_in[11] _6502_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_159_594 VGND VPWR sky130_fd_sc_hd__decap_12
X_3714_ _3711_/A _3759_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_174_520 VGND VPWR sky130_fd_sc_hd__decap_12
X_4694_ _4678_/X _4682_/X _4678_/X _4682_/X _4694_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7482_ _7482_/HI la_data_out[9] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_147_756 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_609 VGND VPWR sky130_fd_sc_hd__fill_1
X_6433_ _6408_/A _6408_/B _6408_/X _6432_/X _6433_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_162_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_597 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_288 VGND VPWR sky130_fd_sc_hd__decap_12
X_6364_ wbs_dat_i[5] _6364_/B _6364_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_115_631 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_269 VGND VPWR sky130_fd_sc_hd__decap_12
X_5315_ _4756_/X _4760_/X _4756_/X _4760_/X _5315_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_141 VGND VPWR sky130_fd_sc_hd__decap_12
X_6295_ _6211_/A _6295_/B _7752_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_170_770 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_472 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_612 VGND VPWR sky130_fd_sc_hd__decap_4
X_5246_ _5232_/X _5236_/X _5235_/X _5246_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_64_1171 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_762 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1144 VGND VPWR sky130_fd_sc_hd__decap_12
X_5177_ _4743_/A _3930_/A _5177_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_96_570 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_581 VGND VPWR sky130_fd_sc_hd__decap_6
X_4128_ _4127_/A _4127_/B _4127_/X _4128_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_83_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_968 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_776 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_15 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_927 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_309 VGND VPWR sky130_fd_sc_hd__decap_12
X_4059_ _4059_/A _4059_/B _4059_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_71_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_459 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_304 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_315 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_623 VGND VPWR sky130_fd_sc_hd__decap_6
X_7818_ _7404_/Y _3914_/A _7810_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_326 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_337 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_645 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_348 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_359 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_818 VGND VPWR sky130_fd_sc_hd__decap_12
X_7749_ _7749_/D _7749_/Q _7746_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_178_870 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_879 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1126 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_767 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_428 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_491 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1041 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_1090 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_623 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_1085 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_931 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_986 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_570 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1214 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_716 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_456 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_916 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_927 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_169 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_724 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_651 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_386 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1056 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_476 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_306 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_380 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_745 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_570 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_907 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_406 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1051 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1013 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_984 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_910 VGND VPWR sky130_fd_sc_hd__decap_12
X_5100_ _5162_/A _4830_/B _5100_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_174_1174 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_780 VGND VPWR sky130_fd_sc_hd__decap_12
X_6080_ _6081_/A _6079_/X _6080_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_32_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1027 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_291 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_965 VGND VPWR sky130_fd_sc_hd__fill_1
X_5031_ _5016_/X _5029_/X _5030_/Y _5032_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_97_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_902 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_710 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1024 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_434 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_968 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_1079 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_573 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_629 VGND VPWR sky130_fd_sc_hd__decap_12
X_6982_ _6941_/Y _6942_/Y _6981_/X _6982_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_93_595 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1240 VGND VPWR sky130_fd_sc_hd__fill_1
X_5933_ _5787_/A _4488_/Y _5933_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_111_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_779 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1270 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_623 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1179 VGND VPWR sky130_fd_sc_hd__decap_12
X_5864_ _4742_/A _5835_/B _5864_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_21_301 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_1276 VGND VPWR sky130_fd_sc_hd__fill_1
X_7603_ _7246_/X _7181_/A _7729_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_167_818 VGND VPWR sky130_fd_sc_hd__decap_3
X_4815_ _4814_/A _4814_/B _4891_/B _4815_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_178_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_947 VGND VPWR sky130_fd_sc_hd__decap_12
X_5795_ _5792_/X _5793_/X _5794_/X _5795_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_166_328 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_367 VGND VPWR sky130_fd_sc_hd__decap_12
X_7534_ _7534_/HI la_data_out[61] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_147_520 VGND VPWR sky130_fd_sc_hd__decap_12
X_4746_ _4741_/X _4745_/X _4744_/X _4746_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_175_840 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_918 VGND VPWR sky130_fd_sc_hd__fill_1
X_7465_ _7465_/HI io_out[30] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_147_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_4677_ _4665_/X _4669_/X _4665_/X _4669_/X _4677_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_147_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1074 VGND VPWR sky130_fd_sc_hd__decap_12
X_6416_ la_data_in[115] _6417_/B VGND VPWR sky130_fd_sc_hd__inv_8
X_7396_ io_in[35] _7396_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_89_802 VGND VPWR sky130_fd_sc_hd__fill_2
X_6347_ _6350_/A _6347_/B _6347_/C _6347_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_192_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_932 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_216 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_868 VGND VPWR sky130_fd_sc_hd__decap_12
X_6278_ _6219_/X _6276_/X _6277_/Y _7756_/D VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_131_965 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_678 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1269 VGND VPWR sky130_fd_sc_hd__decap_8
X_5229_ _5224_/X _5225_/X _5224_/X _5225_/X _5229_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_102_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_708 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1007 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_919 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_101 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_150 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_684 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_134 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_68 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_145 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_806 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_156 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_464 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_167 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_654 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_178 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_879 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_189 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_648 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_969 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_890 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1095 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_1210 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_500 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_748 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_1008 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_83 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_544 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_887 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_729 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_386 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_494 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_0_wb_clk_i clkbuf_1_1_1_wb_clk_i/X clkbuf_2_3_0_wb_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_97_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_367 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_987 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1085 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1077 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_510 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_724 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_426 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1265 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_297 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_543 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_779 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_919 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_932 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_651 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_971 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_418 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_442 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_818 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_497 VGND VPWR sky130_fd_sc_hd__decap_12
X_4600_ _4595_/X _4599_/X _4595_/X _4599_/X _4600_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5580_ _5580_/A _5581_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_175_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1023 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_607 VGND VPWR sky130_fd_sc_hd__decap_3
X_4531_ _7730_/Q _4532_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_129_575 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1187 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_1203 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_681 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_883 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_74 VGND VPWR sky130_fd_sc_hd__decap_12
X_7250_ wbs_stb_i _3695_/A wbs_ack_o VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_176_1225 VGND VPWR sky130_fd_sc_hd__decap_12
X_4462_ _4462_/A _4462_/B _4462_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_171_342 VGND VPWR sky130_fd_sc_hd__decap_12
X_6201_ _5565_/X _6201_/B _6202_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_172_898 VGND VPWR sky130_fd_sc_hd__decap_12
X_4393_ _5130_/A _4647_/B _4393_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7181_ _7181_/A _7181_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_6132_ _4317_/X _6125_/X _6132_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_98_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_965 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_762 VGND VPWR sky130_fd_sc_hd__fill_1
X_6063_ _6033_/A _6061_/X _6311_/B _6063_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_85_315 VGND VPWR sky130_fd_sc_hd__decap_8
X_5014_ _6018_/A _6018_/B _5014_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_85_359 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1237 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_245 VGND VPWR sky130_fd_sc_hd__decap_12
X_6965_ _6965_/A _6965_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_3619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_960 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1070 VGND VPWR sky130_fd_sc_hd__decap_12
X_5916_ _5914_/X _5915_/X _5916_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_2918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6896_ _6876_/X _6894_/X _6895_/Y _6896_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XPHY_2929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1013 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_306 VGND VPWR sky130_fd_sc_hd__decap_12
X_5847_ _5843_/X _5844_/X _5845_/Y _5846_/X _5847_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_22_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_946 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_339 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_968 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_849 VGND VPWR sky130_fd_sc_hd__decap_12
X_5778_ _5776_/X _5777_/X _5778_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7517_ _7517_/HI la_data_out[44] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_182_629 VGND VPWR sky130_fd_sc_hd__decap_12
X_4729_ _4713_/X _4727_/X _4713_/X _4727_/X _4729_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_120_1268 VGND VPWR sky130_fd_sc_hd__decap_8
X_7448_ _7448_/HI io_out[13] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_174_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_876 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_707 VGND VPWR sky130_fd_sc_hd__decap_12
X_7379_ _4540_/Y _7354_/X _7378_/X wbs_dat_o[22] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_150_548 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_805 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_698 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_819 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_231 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_404 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_938 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_370 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_4810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1012 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_993 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1192 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1154 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1162 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_733 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_626 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_102 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_895 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_567 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_330 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_504 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_684 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1128 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_646 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1188 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_348 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_321 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_855 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_573 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_212 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_392 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_245 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_1252 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_1210 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1274 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_587 VGND VPWR sky130_fd_sc_hd__decap_12
X_6750_ _7666_/Q la_data_in[32] _6814_/A VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_50_215 VGND VPWR sky130_fd_sc_hd__decap_6
X_3962_ _3913_/Y _3961_/X _3962_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_91_1123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_395 VGND VPWR sky130_fd_sc_hd__fill_2
X_5701_ _5627_/X _5628_/X _5627_/X _5628_/X _5701_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6681_ _6656_/X _6679_/X _6680_/Y _6681_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_56_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_440 VGND VPWR sky130_fd_sc_hd__decap_6
X_3893_ _3892_/Y _5787_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_176_434 VGND VPWR sky130_fd_sc_hd__decap_12
X_5632_ _5632_/A _5632_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_177_968 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_495 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_467 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_618 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_309 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_501 VGND VPWR sky130_fd_sc_hd__decap_12
X_5563_ _5551_/X _5560_/X _5561_/X _5562_/X _5564_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_145_821 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_437 VGND VPWR sky130_fd_sc_hd__decap_12
X_7302_ _5867_/A _7280_/X _7298_/X _7301_/Y wbs_dat_o[6] VGND VPWR sky130_fd_sc_hd__a211o_4
X_4514_ _4514_/A _4570_/B _4514_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_5494_ _5479_/X _5485_/X _5492_/X _5493_/X _5494_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_172_662 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_353 VGND VPWR sky130_fd_sc_hd__decap_12
X_7233_ _7192_/X _7231_/X _7232_/Y _7233_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_137_1006 VGND VPWR sky130_fd_sc_hd__decap_12
X_4445_ _4322_/Y _4384_/Y _4445_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_104_239 VGND VPWR sky130_fd_sc_hd__decap_12
X_7164_ la_data_in[103] _7165_/B VGND VPWR sky130_fd_sc_hd__inv_8
X_4376_ _7777_/Q _4376_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_99_974 VGND VPWR sky130_fd_sc_hd__fill_2
X_6115_ _6112_/Y _6113_/X _6116_/C VGND VPWR sky130_fd_sc_hd__and2_4
X_7095_ _7095_/A _7095_/B _7095_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_140_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_412 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1130 VGND VPWR sky130_fd_sc_hd__decap_12
X_6046_ _7348_/A _6050_/B _6045_/Y _7793_/D VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_100_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_1050 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_562 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1094 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_4128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1029 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_727 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6948_ la_data_in[71] _6949_/B VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_2704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_790 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_59 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_440 VGND VPWR sky130_fd_sc_hd__decap_12
X_6879_ _6822_/Y _6824_/B _6824_/X _6878_/X _6880_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XPHY_2759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_412 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_905 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1062 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_876 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_1253 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_898 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_559 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_889 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_107 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1044 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_724 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_1172 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_392 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1099 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_82 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_4640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_215 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_379 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_570 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_259 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_440 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_581 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_579 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_1107 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_968 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_938 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_466 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_426 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1184 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1203 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_386 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1217 VGND VPWR sky130_fd_sc_hd__decap_3
X_4230_ _4227_/X _4229_/X _4240_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_141_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1091 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_922 VGND VPWR sky130_fd_sc_hd__decap_12
X_4161_ _4505_/A _4218_/B _4161_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_122_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_123 VGND VPWR sky130_fd_sc_hd__decap_12
X_4092_ _4092_/A _4091_/X _4092_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_96_999 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1223 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_502 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_727 VGND VPWR sky130_fd_sc_hd__decap_3
X_6802_ _6738_/X _6758_/B _6802_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_7782_ _7782_/D _4070_/A _7746_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_24_749 VGND VPWR sky130_fd_sc_hd__decap_12
X_4994_ _4415_/X _4416_/X _4415_/X _4416_/X _4994_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_196_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_1093 VGND VPWR sky130_fd_sc_hd__decap_4
X_6733_ _7672_/Q _6735_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_205_891 VGND VPWR sky130_fd_sc_hd__decap_12
X_3945_ _4189_/A _3933_/X _3946_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_143_1010 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1013 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_771 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_922 VGND VPWR sky130_fd_sc_hd__decap_12
X_6664_ la_data_in[31] _6663_/Y _6666_/B VGND VPWR sky130_fd_sc_hd__nor2_4
X_3876_ _3875_/Y _3877_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_177_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1065 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_966 VGND VPWR sky130_fd_sc_hd__decap_12
X_5615_ _5072_/A _4612_/B _5615_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_149_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_117 VGND VPWR sky130_fd_sc_hd__decap_12
X_6595_ _6595_/A _6668_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_178_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1224 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_320 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_459 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_768 VGND VPWR sky130_fd_sc_hd__fill_1
X_5546_ _4803_/X _4804_/X _4803_/X _4804_/X _5546_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_145_662 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_684 VGND VPWR sky130_fd_sc_hd__decap_6
X_5477_ _5471_/X _5476_/X _5471_/X _5476_/X _5477_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_155_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_846 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_548 VGND VPWR sky130_fd_sc_hd__fill_1
X_7216_ _7200_/X _7215_/X _7212_/X _7216_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_160_654 VGND VPWR sky130_fd_sc_hd__decap_12
X_4428_ _4898_/A _4512_/B _4428_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_133_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_602 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1153 VGND VPWR sky130_fd_sc_hd__decap_12
X_7147_ _7145_/Y _7147_/B _7147_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_4359_ _4359_/A _4358_/X _4359_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_115_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_27 VGND VPWR sky130_fd_sc_hd__decap_12
X_7078_ _7073_/Y _7074_/Y _7139_/B _7078_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_74_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1224 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_178 VGND VPWR sky130_fd_sc_hd__decap_12
X_6029_ _7327_/A _3967_/X _6060_/A _6029_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_55_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_159 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_800 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_806 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_373 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_215 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_749 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_367 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_877 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1102 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_579 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1162 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1132 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_850 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_220 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_68 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_776 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_724 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_68 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_62 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_746 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_876 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_353 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_159_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_790 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1220 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_697 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1245 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_819 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_1267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1095 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_4470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_855 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_719 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1062 VGND VPWR sky130_fd_sc_hd__decap_12
X_3730_ _4494_/A _4793_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_60_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_793 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_590 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_281 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_618 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_285 VGND VPWR sky130_fd_sc_hd__decap_12
X_5400_ _5378_/X _5379_/X _5378_/X _5379_/X _5400_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_173_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_459 VGND VPWR sky130_fd_sc_hd__decap_12
X_6380_ wbs_dat_i[0] _6334_/B _6381_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_62_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_802 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_971 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_1082 VGND VPWR sky130_fd_sc_hd__decap_12
X_5331_ _5289_/X _5330_/X _5289_/X _5330_/X _5331_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1033 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1044 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1003 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_654 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_345 VGND VPWR sky130_fd_sc_hd__decap_12
X_5262_ _5259_/X _5260_/X _5261_/X _5262_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_173_1036 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_665 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1167 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_900 VGND VPWR sky130_fd_sc_hd__decap_12
X_7001_ _6984_/X _6998_/X _7000_/Y _7646_/D VGND VPWR sky130_fd_sc_hd__o21a_4
X_4213_ _4194_/X _4195_/X _4194_/X _4195_/X _4213_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_5193_ _5184_/X _5190_/X _5191_/X _5192_/X _5193_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_96_730 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_944 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1228 VGND VPWR sky130_fd_sc_hd__decap_12
X_4144_ _4843_/A _4145_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_68_454 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_796 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1111 VGND VPWR sky130_fd_sc_hd__decap_8
X_4075_ _5058_/A _3924_/X _4075_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_37_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1015 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_373 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_395 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_855 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_192 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_7765_ _7765_/D _5292_/A _7769_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_51_365 VGND VPWR sky130_fd_sc_hd__fill_1
X_4977_ _4953_/X _4976_/X _4953_/X _4976_/X _4977_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_337 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_220 VGND VPWR sky130_fd_sc_hd__decap_12
X_6716_ la_data_in[44] _6717_/B VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3928_ _3928_/A _4654_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_211_168 VGND VPWR sky130_fd_sc_hd__decap_12
X_7696_ _6668_/X _6600_/A _7696_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_177_562 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_752 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_938 VGND VPWR sky130_fd_sc_hd__decap_8
X_6647_ _6647_/A _6647_/B _6698_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_50_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_3859_ _3858_/Y _4697_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_192_532 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_297 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_640 VGND VPWR sky130_fd_sc_hd__fill_1
X_6578_ _6586_/A _6545_/X _6578_/C _6578_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_121_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_727 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_929 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_993 VGND VPWR sky130_fd_sc_hd__decap_12
X_5529_ _5525_/X _5528_/X _5525_/X _5528_/X _5529_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_69_1253 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_428 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_1234 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_963 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1128 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_356 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_849 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_909 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_627 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_284 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_126 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1213 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_107 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_74 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_855 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_1219 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1249 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_669 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1090 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_549 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_916 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_404 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_190 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_745 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_245 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1009 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_587 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1274 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1069 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_930 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_82 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_996 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_849 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1053 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1097 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_65 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_76 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_87 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_788 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_980 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_964 VGND VPWR sky130_fd_sc_hd__decap_12
X_4900_ _4897_/X _4900_/B _4900_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_52_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_693 VGND VPWR sky130_fd_sc_hd__decap_8
X_5880_ _5874_/X _5875_/X _5869_/X _5876_/X _5880_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_209_1135 VGND VPWR sky130_fd_sc_hd__fill_1
X_4831_ _4829_/X _4830_/X _4831_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_33_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1168 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1130 VGND VPWR sky130_fd_sc_hd__decap_12
X_7550_ _7550_/HI la_data_out[77] VGND VPWR sky130_fd_sc_hd__conb_1
X_4762_ _4747_/X _4751_/X _4750_/X _4762_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_92_1081 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_318 VGND VPWR sky130_fd_sc_hd__decap_12
X_6501_ _6501_/A _6503_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_3713_ _3693_/X _3712_/X _3717_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_186_370 VGND VPWR sky130_fd_sc_hd__decap_12
X_7481_ _7481_/HI la_data_out[8] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_119_426 VGND VPWR sky130_fd_sc_hd__fill_1
X_4693_ _4684_/X _4685_/X _4684_/X _4685_/X _4693_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_174_532 VGND VPWR sky130_fd_sc_hd__decap_12
X_6432_ _6409_/Y _6410_/Y _6476_/B _6432_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_147_768 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1245 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_1128 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_727 VGND VPWR sky130_fd_sc_hd__decap_12
X_6363_ _6345_/A _6364_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_162_749 VGND VPWR sky130_fd_sc_hd__decap_12
X_5314_ _5161_/X _5165_/X _5164_/X _5314_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_6294_ _5983_/X _6219_/A _6293_/Y _5867_/A _6084_/X _6295_/B VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_102_304 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_793 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_484 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_624 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_698 VGND VPWR sky130_fd_sc_hd__decap_12
X_5245_ _5240_/X _5244_/X _5243_/X _5245_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_102_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1206 VGND VPWR sky130_fd_sc_hd__decap_12
X_5176_ _5176_/A _3938_/A _5176_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_190_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1156 VGND VPWR sky130_fd_sc_hd__decap_3
X_4127_ _4127_/A _4127_/B _4127_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_112_1126 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_608 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1227 VGND VPWR sky130_fd_sc_hd__decap_12
X_4058_ _4583_/A _4126_/B _4059_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_72_939 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_855 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_305 VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_5_0_wb_clk_i clkbuf_2_2_1_wb_clk_i/X clkbuf_3_5_0_wb_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_316 VGND VPWR sky130_fd_sc_hd__decap_3
X_7817_ _7817_/D _3689_/A _7810_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_327 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_983 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_674 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_338 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_825 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_349 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_657 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_836 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_184 VGND VPWR sky130_fd_sc_hd__decap_12
X_7748_ _6312_/X _5946_/A _7746_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_123_1200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_882 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1233 VGND VPWR sky130_fd_sc_hd__decap_12
X_7679_ _6780_/X _7679_/Q _7658_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_177_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_726 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1020 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_963 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_921 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_1097 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1250 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_943 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_240 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1234 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_871 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_728 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_703 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_35_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_939 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_736 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1013 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_663 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_877 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_978 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1038 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_398 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_346 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_713 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_392 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_757 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_513 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_738 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_395 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1063 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_771 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_825 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_1025 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_922 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_996 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_613 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_484 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_847 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1186 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1039 VGND VPWR sky130_fd_sc_hd__decap_8
X_5030_ _5016_/X _5029_/X _5030_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_97_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_722 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1036 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_593 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_958 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_755 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_703 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_468 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_479 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1020 VGND VPWR sky130_fd_sc_hd__decap_8
X_6981_ _7008_/A _7008_/B _6981_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_93_585 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_32 VGND VPWR sky130_fd_sc_hd__decap_12
X_5932_ _3901_/X _4475_/Y _5932_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_20_1086 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_961 VGND VPWR sky130_fd_sc_hd__decap_12
X_5863_ _5860_/X _5861_/X _5862_/X _5863_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_55_1127 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_825 VGND VPWR sky130_fd_sc_hd__decap_12
X_7602_ _7602_/D _7602_/Q _7729_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_179_668 VGND VPWR sky130_fd_sc_hd__decap_3
X_4814_ _4814_/A _4814_/B _4891_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_33_184 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_605 VGND VPWR sky130_fd_sc_hd__decap_12
X_5794_ _5792_/X _5793_/X _5794_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_178_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_959 VGND VPWR sky130_fd_sc_hd__decap_12
X_7533_ _7533_/HI la_data_out[60] VGND VPWR sky130_fd_sc_hd__conb_1
X_4745_ _4742_/X _4743_/X _4744_/X _4745_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_21_379 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_147_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_852 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_245 VGND VPWR sky130_fd_sc_hd__decap_12
X_7464_ _7464_/HI io_out[29] VGND VPWR sky130_fd_sc_hd__conb_1
X_4676_ _4671_/X _4672_/X _4671_/X _4672_/X _4676_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_190_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_1160 VGND VPWR sky130_fd_sc_hd__decap_12
X_6415_ _7717_/Q _6415_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_147_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_7395_ _7394_/Y _7387_/X _7774_/Q _7388_/X wbs_dat_o[28] VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_179_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_440 VGND VPWR sky130_fd_sc_hd__decap_12
X_6346_ wbs_dat_i[10] _6349_/B _6347_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_1_707 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_718 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_410 VGND VPWR sky130_fd_sc_hd__decap_12
X_6277_ _5754_/A _6106_/X _6595_/A _6277_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_163_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_668 VGND VPWR sky130_fd_sc_hd__decap_3
X_5228_ _5120_/X _5227_/X _5120_/X _5227_/X _5228_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_130_487 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1010 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_413 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1081 VGND VPWR sky130_fd_sc_hd__decap_12
X_5159_ _5156_/X _5157_/X _5158_/X _5159_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_57_788 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_922 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_257 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_102 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_663 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_113 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_123 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_135 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_791 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_146 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_476 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_168 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_318 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_179 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_666 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_1060 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_512 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_1159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_579 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_440 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_398 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_806 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_999 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_773 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1097 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_574 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_788 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_1067 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_1127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_287 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_555 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_410 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_663 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_983 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_764 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_786 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_307 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_80 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1171 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_830 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1035 VGND VPWR sky130_fd_sc_hd__decap_12
X_4530_ _4530_/A _4495_/X _4530_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_7_31 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_587 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_1245 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_693 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_4461_ _4461_/A _4461_/B _4462_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_7_86 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_1237 VGND VPWR sky130_fd_sc_hd__decap_12
X_6200_ _5583_/X _6199_/X _6004_/B _6201_/B VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_171_354 VGND VPWR sky130_fd_sc_hd__decap_12
X_7180_ _7180_/A _7180_/B _7180_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_144_579 VGND VPWR sky130_fd_sc_hd__fill_1
X_4392_ _5052_/A _4653_/B _4392_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_113_911 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_600 VGND VPWR sky130_fd_sc_hd__decap_8
X_6131_ _6128_/X _6129_/Y _6130_/X _7781_/D VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_112_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_977 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_508 VGND VPWR sky130_fd_sc_hd__decap_8
X_6062_ _6139_/A _6311_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_26_1240 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1210 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_891 VGND VPWR sky130_fd_sc_hd__fill_2
X_5013_ _5013_/A _6018_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_39_733 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_861 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_872 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_1249 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_747 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6964_ _6962_/Y _6963_/Y _6964_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_53_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_972 VGND VPWR sky130_fd_sc_hd__decap_4
X_5915_ _3900_/Y _4480_/Y _5915_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_2908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6895_ _6876_/X _6894_/X _6811_/X _6895_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XPHY_2919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1030 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1082 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_471 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_482 VGND VPWR sky130_fd_sc_hd__decap_12
X_5846_ _5843_/X _5844_/X _5843_/X _5844_/X _5846_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_195_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_318 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_649 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_767 VGND VPWR sky130_fd_sc_hd__decap_12
X_5777_ _5664_/X _5675_/X _5643_/X _5676_/X _5777_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_194_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1203 VGND VPWR sky130_fd_sc_hd__decap_12
X_4728_ _4526_/X _4527_/X _4526_/X _4527_/X _4728_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7516_ _7516_/HI la_data_out[43] VGND VPWR sky130_fd_sc_hd__conb_1
X_7447_ _7447_/HI io_out[12] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_163_844 VGND VPWR sky130_fd_sc_hd__decap_8
X_4659_ _4655_/X _4657_/X _4658_/X _4659_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_163_855 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_888 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_719 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_900 VGND VPWR sky130_fd_sc_hd__decap_12
X_7378_ _4539_/A _7370_/X _7377_/Y _7364_/X _7378_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_162_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1110 VGND VPWR sky130_fd_sc_hd__decap_12
X_6329_ _6332_/A _6329_/B _6329_/C _6329_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_27_1004 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_1012 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_741 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_1045 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_817 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_574 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_416 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_511 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1130 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1103 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1136 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_638 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_186_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_114 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1013 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_811 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_663 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_516 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1178 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_947 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_958 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_338 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_658 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_541 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_883 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_360 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_257 VGND VPWR sky130_fd_sc_hd__decap_12
X_3961_ _3918_/X _3924_/X _3961_/C _3961_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_56_1222 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_509 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_599 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_471 VGND VPWR sky130_fd_sc_hd__decap_3
X_5700_ _5696_/X _5699_/X _5700_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_182_1241 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_774 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1135 VGND VPWR sky130_fd_sc_hd__decap_8
X_6680_ _6656_/X _6679_/X _6670_/X _6680_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_188_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1217 VGND VPWR sky130_fd_sc_hd__decap_3
X_3892_ _7795_/Q _3892_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_52_1108 VGND VPWR sky130_fd_sc_hd__fill_1
X_5631_ _5597_/X _5613_/X _5629_/X _5630_/X _5631_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_176_446 VGND VPWR sky130_fd_sc_hd__decap_12
X_5562_ _5551_/X _5560_/X _5551_/X _5560_/X _5562_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_117_513 VGND VPWR sky130_fd_sc_hd__decap_12
X_7301_ _5137_/A _7293_/X _7300_/X _7301_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_145_833 VGND VPWR sky130_fd_sc_hd__decap_12
X_4513_ _4513_/A _4569_/B _4515_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_191_449 VGND VPWR sky130_fd_sc_hd__decap_12
X_5493_ _5479_/X _5485_/X _5479_/X _5485_/X _5493_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_145_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_557 VGND VPWR sky130_fd_sc_hd__decap_12
X_7232_ _7192_/X _7231_/X _6085_/X _7232_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_4444_ _4443_/X _4444_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_144_365 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1067 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_1018 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1078 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_398 VGND VPWR sky130_fd_sc_hd__decap_12
X_7163_ _7609_/Q _7163_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4375_ _4325_/X _4353_/X _4373_/X _4374_/X _4375_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_6114_ _6112_/Y _6113_/X _6114_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_98_463 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_914 VGND VPWR sky130_fd_sc_hd__fill_1
X_7094_ _7037_/Y _7038_/Y _7039_/X _7093_/X _7095_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_140_593 VGND VPWR sky130_fd_sc_hd__decap_8
X_6045_ _7348_/A _6050_/B _6595_/A _6045_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_58_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_202 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_566 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_352 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_419 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1038 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_279 VGND VPWR sky130_fd_sc_hd__decap_12
X_6947_ _6947_/A _6947_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_2705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_739 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_27 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6878_ _6825_/Y _6827_/B _6827_/X _6877_/X _6878_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_50_750 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_452 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_424 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_195_733 VGND VPWR sky130_fd_sc_hd__decap_3
X_5829_ _5827_/X _5828_/X _5829_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_139_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_928 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_788 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1191 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_471 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_1107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_482 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_538 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_345 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_356 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_284 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1181 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_190 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_257 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_503 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_227 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_903 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_401 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_1119 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_478 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_489 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_693 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_1242 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_825 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_847 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_32 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_379 VGND VPWR sky130_fd_sc_hd__decap_12
X_4160_ _4513_/A _4505_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_96_934 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_135 VGND VPWR sky130_fd_sc_hd__decap_12
X_4091_ _4072_/X _4088_/X _4089_/X _4090_/X _4091_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_23_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_675 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1235 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1268 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_672 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_886 VGND VPWR sky130_fd_sc_hd__decap_12
X_6801_ _6759_/X _6799_/X _6800_/Y _6801_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_208_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_514 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_683 VGND VPWR sky130_fd_sc_hd__decap_12
X_4993_ _4431_/X _4432_/X _4431_/X _4432_/X _4993_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7781_ _7781_/D _7781_/Q _7746_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_23_216 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1030 VGND VPWR sky130_fd_sc_hd__fill_2
X_3944_ _3693_/X _3924_/X _3946_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_6732_ _6730_/Y _6732_/B _6732_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_32_761 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_1022 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1025 VGND VPWR sky130_fd_sc_hd__decap_12
X_6663_ io_out[1] _6663_/B _6663_/Y VGND VPWR sky130_fd_sc_hd__xnor2_4
XFILLER_32_783 VGND VPWR sky130_fd_sc_hd__decap_12
X_3875_ _3875_/A _3875_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_20_934 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_703 VGND VPWR sky130_fd_sc_hd__decap_12
X_5614_ _5606_/X _5610_/X _5606_/X _5610_/X _5614_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_177_788 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1077 VGND VPWR sky130_fd_sc_hd__decap_6
X_6594_ _6536_/X _6592_/X _6593_/Y _7700_/D VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_176_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_978 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_833 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_449 VGND VPWR sky130_fd_sc_hd__decap_8
X_5545_ _5521_/X _5542_/X _5543_/X _5544_/X _5548_/A VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_30_1236 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_332 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_877 VGND VPWR sky130_fd_sc_hd__decap_8
X_5476_ _5474_/X _5475_/X _5474_/X _5475_/X _5476_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_172_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_516 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_324 VGND VPWR sky130_fd_sc_hd__decap_12
X_4427_ _4612_/B _4512_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_7215_ _7614_/Q la_data_in[108] _7150_/X _7215_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_160_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1192 VGND VPWR sky130_fd_sc_hd__decap_12
X_7146_ la_data_in[109] _7147_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_63_1034 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_1215 VGND VPWR sky130_fd_sc_hd__decap_12
X_4358_ _3720_/A _4505_/B _4358_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_48_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_794 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1165 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1198 VGND VPWR sky130_fd_sc_hd__decap_12
X_7077_ _7077_/A _7138_/B _7139_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_171_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_809 VGND VPWR sky130_fd_sc_hd__decap_12
X_4289_ _4289_/A _4289_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_189_1236 VGND VPWR sky130_fd_sc_hd__decap_12
X_6028_ _6028_/A _6028_/B _6027_/Y _6060_/A VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_86_488 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_500 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_190 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_3203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_385 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_227 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_508 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_32 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1130 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_379 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1114 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1174 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1144 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_862 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_794 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_350 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_361 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_916 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_202 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_949 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_758 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_888 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_460 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1062 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_666 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_145_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_508 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1123 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_1145 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_444 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_135 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_197 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_650 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1063 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_678 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_322 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_867 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_344 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1252 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_3770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_722 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_891 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1274 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1074 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_928 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_253 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_630 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_297 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_80 VGND VPWR sky130_fd_sc_hd__decap_12
X_5330_ _5328_/X _5329_/X _5328_/X _5329_/X _5330_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_115_814 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_960 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1094 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_696 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_324 VGND VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_7_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/A _7769_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_177_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1067 VGND VPWR sky130_fd_sc_hd__fill_1
X_5261_ _5259_/X _5260_/X _5261_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_114_357 VGND VPWR sky130_fd_sc_hd__decap_12
X_7000_ _6984_/X _6998_/X _6999_/X _7000_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_142_677 VGND VPWR sky130_fd_sc_hd__decap_12
X_4212_ _4197_/Y _4198_/X _4197_/Y _4198_/X _4251_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_87_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_912 VGND VPWR sky130_fd_sc_hd__decap_3
X_5192_ _5184_/X _5190_/X _5184_/X _5190_/X _5192_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_69_956 VGND VPWR sky130_fd_sc_hd__decap_12
X_4143_ _4143_/A _4843_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_96_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1270 VGND VPWR sky130_fd_sc_hd__decap_6
X_4074_ _5069_/A _3933_/X _4074_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_205_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_959 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1062 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1032 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_300 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_1087 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1027 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_806 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_867 VGND VPWR sky130_fd_sc_hd__decap_12
X_7764_ _7764_/D _5062_/A _7769_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_211_125 VGND VPWR sky130_fd_sc_hd__decap_12
X_4976_ _4974_/X _4975_/X _4974_/X _4975_/X _4976_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_208 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_349 VGND VPWR sky130_fd_sc_hd__decap_12
X_6715_ _6715_/A _6717_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_3927_ _3718_/A _3919_/A _3927_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_177_541 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_232 VGND VPWR sky130_fd_sc_hd__decap_12
X_7695_ _6672_/X _7695_/Q _7758_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_3858_ _3858_/A _3858_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_6646_ _6635_/A _6634_/Y _6635_/X _6645_/X _6647_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_164_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1180 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1191 VGND VPWR sky130_fd_sc_hd__decap_12
X_3789_ _4459_/A _3767_/B _3791_/B VGND VPWR sky130_fd_sc_hd__and2_4
X_6577_ _6545_/A _6544_/X _6578_/C VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_69_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1172 VGND VPWR sky130_fd_sc_hd__decap_12
X_5528_ _5526_/X _5527_/X _5526_/X _5527_/X _5528_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_133_611 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1276 VGND VPWR sky130_fd_sc_hd__fill_1
X_5459_ _6006_/A _6006_/B _5459_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_156_1246 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_709 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_452 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_580 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_349 VGND VPWR sky130_fd_sc_hd__decap_12
X_7129_ _7066_/X _7081_/B _7129_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_8_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_541 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_138 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1099 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_801 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_886 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_199_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1225 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_672 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_182 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_839 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_867 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_558 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_569 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_517 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_528 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_906 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_552 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_928 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_223 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_641 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_268 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_599 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_685 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_780 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_791 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_942 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_891 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_1062 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_764 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1065 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_11 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_831 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_992 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_480 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_396 VGND VPWR sky130_fd_sc_hd__fill_1
X_4830_ _4485_/A _4830_/B _4830_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_209_1158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_141 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1180 VGND VPWR sky130_fd_sc_hd__fill_2
X_4761_ _4756_/X _4760_/X _4759_/X _4761_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_57_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_541 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_703 VGND VPWR sky130_fd_sc_hd__decap_12
X_3712_ _3757_/A _3712_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_6500_ _6500_/A _6500_/B _6500_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_174_500 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1003 VGND VPWR sky130_fd_sc_hd__decap_4
X_7480_ _7480_/HI la_data_out[7] VGND VPWR sky130_fd_sc_hd__conb_1
X_4692_ _4687_/X _4688_/X _4687_/X _4688_/X _4692_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_382 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_544 VGND VPWR sky130_fd_sc_hd__decap_12
X_6431_ _6431_/A _6431_/B _6476_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_140_1069 VGND VPWR sky130_fd_sc_hd__decap_12
X_6362_ _4299_/X _6373_/B _6365_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_162_739 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_611 VGND VPWR sky130_fd_sc_hd__decap_12
X_5313_ _5299_/X _5312_/X _5299_/X _5312_/X _5313_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_115_644 VGND VPWR sky130_fd_sc_hd__decap_8
X_6293_ _5983_/A _6293_/B _6293_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_170_750 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_655 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_154 VGND VPWR sky130_fd_sc_hd__decap_12
X_5244_ _5241_/X _5242_/X _5243_/X _5244_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_102_316 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_496 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_636 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_349 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_1170 VGND VPWR sky130_fd_sc_hd__decap_12
X_5175_ _4741_/X _4745_/X _4741_/X _4745_/X _5175_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_116_1252 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_1214 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_263 VGND VPWR sky130_fd_sc_hd__decap_12
X_4126_ _4539_/A _4126_/B _4127_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_69_797 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1176 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_1059 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_425 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_594 VGND VPWR sky130_fd_sc_hd__decap_12
X_4057_ _4923_/B _4126_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_186_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_672 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_642 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_306 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1072 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_867 VGND VPWR sky130_fd_sc_hd__decap_12
X_7816_ _3725_/Y _3718_/A _7810_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_149_1083 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_317 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_328 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_339 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_27 VGND VPWR sky130_fd_sc_hd__decap_8
X_7747_ _7747_/D _7747_/Q _7746_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_71_1122 VGND VPWR sky130_fd_sc_hd__decap_12
X_4959_ _4959_/A _4959_/B _4959_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_200_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1212 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1106 VGND VPWR sky130_fd_sc_hd__decap_12
X_7678_ _6783_/X _6715_/A _7658_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_123_1245 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1177 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_533 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_842 VGND VPWR sky130_fd_sc_hd__decap_12
X_6629_ _6627_/Y _6628_/Y _6627_/Y _6628_/Y _6695_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_180_503 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_471 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_193_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_622 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_791 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1062 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_900 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_794 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_955 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1246 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_883 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_745 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_959 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_907 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_469 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_300 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_171 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1150 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_940 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1044 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_193 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1172 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_1025 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_135 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_185 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_489 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1191 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_725 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_202 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_550 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_510 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_532 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_706 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1020 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_1151 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_430 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_174_1121 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_964 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_603 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_783 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1097 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_625 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_314 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_859 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_745 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1048 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_918 VGND VPWR sky130_fd_sc_hd__decap_12
X_6980_ _6944_/Y _6945_/Y _7012_/B _7008_/B VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_111_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_428 VGND VPWR sky130_fd_sc_hd__decap_12
X_5931_ _3877_/A _4532_/A _5931_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_202_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_620 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1253 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1148 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_951 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_642 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_973 VGND VPWR sky130_fd_sc_hd__decap_12
X_5862_ _5860_/X _5861_/X _5862_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_90_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_1139 VGND VPWR sky130_fd_sc_hd__decap_12
X_7601_ _7249_/X _3695_/A _7785_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_22_837 VGND VPWR sky130_fd_sc_hd__decap_6
X_4813_ _4813_/A _4813_/B _4814_/B VGND VPWR sky130_fd_sc_hd__and2_4
X_5793_ _4742_/A _4482_/A _5793_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_166_308 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_617 VGND VPWR sky130_fd_sc_hd__decap_12
X_7532_ _7532_/HI la_data_out[59] VGND VPWR sky130_fd_sc_hd__conb_1
X_4744_ _4742_/X _4743_/X _4744_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_30_870 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_190 VGND VPWR sky130_fd_sc_hd__decap_12
X_4675_ _4638_/X _4674_/X _4638_/X _4674_/X _4675_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7463_ _7463_/HI io_out[28] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_119_257 VGND VPWR sky130_fd_sc_hd__decap_12
X_6414_ _6412_/Y _6413_/Y _6412_/Y _6413_/Y _6429_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_1172 VGND VPWR sky130_fd_sc_hd__decap_12
X_7394_ io_in[34] _7394_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_174_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_227 VGND VPWR sky130_fd_sc_hd__decap_12
X_6345_ _6345_/A _6349_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_131_901 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_614 VGND VPWR sky130_fd_sc_hd__decap_12
X_6276_ _5857_/X _5990_/B _5990_/X _6276_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_143_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1219 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_218 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_422 VGND VPWR sky130_fd_sc_hd__decap_12
X_5227_ _5211_/X _5226_/X _5211_/X _5226_/X _5227_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_69_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1184 VGND VPWR sky130_fd_sc_hd__decap_8
X_5158_ _5156_/X _5157_/X _5158_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_29_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_1093 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_391 VGND VPWR sky130_fd_sc_hd__decap_6
X_4109_ _4070_/Y _4095_/X _4070_/Y _4095_/X _4109_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_553 VGND VPWR sky130_fd_sc_hd__decap_12
X_5089_ _5084_/X _5088_/X _5087_/X _5089_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_56_288 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_480 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_934 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_269 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_103 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_1217 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_125 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_826 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_905 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_837 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_136 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_916 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_147 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_812 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_193_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_588 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_986 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1021 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1081 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_211 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1245 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_82 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_93 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_5 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_567 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_675 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_956 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_995 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_617 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_319 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1150 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1183 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_168_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_971 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1047 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_43 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_352 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1126 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_863 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1069 VGND VPWR sky130_fd_sc_hd__decap_12
X_4460_ _4554_/A _4460_/B _4462_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_183_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1249 VGND VPWR sky130_fd_sc_hd__fill_2
X_4391_ _4328_/X _4332_/X _4328_/X _4332_/X _4391_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_194_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_208 VGND VPWR sky130_fd_sc_hd__decap_12
X_6130_ _4150_/Y _6103_/X _6092_/X _6130_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_125_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_422 VGND VPWR sky130_fd_sc_hd__decap_8
X_6061_ _3967_/X _6072_/B _6061_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_140_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_678 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_689 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_701 VGND VPWR sky130_fd_sc_hd__decap_8
X_5012_ _5012_/A _6018_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_100_628 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1274 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_1149 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_597 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1081 VGND VPWR sky130_fd_sc_hd__decap_4
X_6963_ la_data_in[66] _6963_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_183_1209 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_480 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_1050 VGND VPWR sky130_fd_sc_hd__fill_2
X_5914_ _3892_/Y _4475_/Y _5914_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_53_269 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6894_ _7661_/Q la_data_in[59] _6830_/X _6894_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_146_1042 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1094 VGND VPWR sky130_fd_sc_hd__decap_4
X_5845_ _7753_/Q _5845_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_34_494 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1097 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_678 VGND VPWR sky130_fd_sc_hd__decap_12
X_5776_ _5770_/X _5771_/X _5770_/X _5771_/X _5776_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_210_779 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1245 VGND VPWR sky130_fd_sc_hd__decap_12
X_7515_ _7515_/HI la_data_out[42] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_147_330 VGND VPWR sky130_fd_sc_hd__decap_12
X_4727_ _4714_/X _4724_/X _4725_/X _4726_/X _4727_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_120_1215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_672 VGND VPWR sky130_fd_sc_hd__decap_12
X_7446_ _7446_/HI io_out[11] VGND VPWR sky130_fd_sc_hd__conb_1
X_4658_ _4655_/X _4657_/X _4658_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_190_642 VGND VPWR sky130_fd_sc_hd__decap_8
X_7377_ io_in[28] _7377_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4589_ _4589_/A _4546_/B _4589_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_104_912 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1021 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1160 VGND VPWR sky130_fd_sc_hd__decap_12
X_6328_ wbs_dat_i[15] _6338_/B _6329_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_143_580 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1122 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_794 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_934 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1065 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_1193 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1024 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_678 VGND VPWR sky130_fd_sc_hd__fill_1
X_6259_ _6256_/X _6258_/X _6057_/A _6259_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_153_1057 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_829 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_211 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_350 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1172 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_764 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_431 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1189 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_1148 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_627 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_126 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_661 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_1025 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1069 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1020 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_1031 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_528 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1097 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_851 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1160 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_1221 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_940 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_353 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_1097 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_269 VGND VPWR sky130_fd_sc_hd__decap_8
X_3960_ _3926_/X _3958_/X _3959_/Y _3961_/C VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_95_1261 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_375 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_910 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1234 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_764 VGND VPWR sky130_fd_sc_hd__decap_3
X_3891_ _3866_/X _3891_/B _3891_/C _7796_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_182_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_786 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_1215 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_5630_ _5597_/X _5613_/X _5597_/X _5613_/X _5630_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_85_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_330 VGND VPWR sky130_fd_sc_hd__decap_12
X_5561_ _5555_/X _5556_/X _5554_/X _5557_/X _5561_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_106_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_672 VGND VPWR sky130_fd_sc_hd__fill_2
X_7300_ _7299_/Y _7300_/B _7300_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4512_ _4512_/A _4512_/B _4512_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_5492_ _5489_/X _5490_/X _5491_/X _5492_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_145_845 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_170 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_867 VGND VPWR sky130_fd_sc_hd__decap_12
X_7231_ _7608_/Q la_data_in[102] _7168_/X _7231_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_208_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_569 VGND VPWR sky130_fd_sc_hd__decap_12
X_4443_ _4443_/A _4443_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_160_837 VGND VPWR sky130_fd_sc_hd__decap_4
X_4374_ _4325_/X _4353_/X _4325_/X _4353_/X _4374_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7162_ _7160_/Y _7161_/Y _7160_/Y _7161_/Y _7226_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_171_196 VGND VPWR sky130_fd_sc_hd__decap_12
X_6113_ _4208_/X _6096_/X _4202_/X _6113_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_7093_ _7040_/Y _7041_/Y _7042_/X _7092_/X _7093_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_99_998 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_263 VGND VPWR sky130_fd_sc_hd__decap_12
X_6044_ _6044_/A _6595_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_86_648 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_436 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_18 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1030 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_586 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1104 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_556 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_247 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1069 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_578 VGND VPWR sky130_fd_sc_hd__fill_2
X_6946_ _6944_/Y _6945_/Y _6944_/Y _6945_/Y _6946_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_3429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_898 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_206 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_39 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6877_ _6830_/A _6830_/B _6830_/X _6876_/X _6877_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_169_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_510 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_762 VGND VPWR sky130_fd_sc_hd__fill_1
X_5828_ _5787_/A _4361_/Y _5828_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_5759_ _5747_/X _5748_/X _5757_/X _5758_/X _5759_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_120_1001 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_608 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1211 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_480 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_631 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_536 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1067 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_32 VGND VPWR sky130_fd_sc_hd__decap_12
X_7429_ io_oeb[24] _7429_/LO VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_162_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_686 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_826 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_494 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_764 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_786 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_296 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_62 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_849 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_353 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_269 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_515 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_910 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_239 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_948 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_424 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_406 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1191 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_672 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_641 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_604 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_80 VGND VPWR sky130_fd_sc_hd__decap_12
X_4090_ _4083_/X _4086_/X _4090_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_67_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_778 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1203 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_361 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_895 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_687 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1247 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_342 VGND VPWR sky130_fd_sc_hd__decap_12
X_6800_ _6759_/X _6799_/X _6785_/X _6800_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_7780_ _7780_/D _7780_/Q _7746_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_898 VGND VPWR sky130_fd_sc_hd__decap_12
X_4992_ _4437_/X _4438_/X _4437_/X _4438_/X _4992_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_91_695 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_526 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_781 VGND VPWR sky130_fd_sc_hd__decap_12
X_6731_ la_data_in[39] _6732_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_189_550 VGND VPWR sky130_fd_sc_hd__decap_12
X_3943_ _3935_/Y _3942_/X _3934_/X _3943_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_210_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_712 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1001 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_583 VGND VPWR sky130_fd_sc_hd__decap_12
X_6662_ _6600_/Y _6601_/Y _6661_/X _6663_/B VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_143_1034 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_1154 VGND VPWR sky130_fd_sc_hd__decap_12
X_3874_ _3866_/X _3874_/B _3874_/C _7798_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_182_1094 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_795 VGND VPWR sky130_fd_sc_hd__decap_12
X_5613_ _5604_/X _5612_/X _5604_/X _5612_/X _5613_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_137_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_715 VGND VPWR sky130_fd_sc_hd__decap_12
X_6593_ _6536_/X _6592_/X _6572_/X _6593_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_176_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_620 VGND VPWR sky130_fd_sc_hd__decap_12
X_5544_ _5521_/X _5542_/X _5521_/X _5542_/X _5544_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_129_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_940 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_1248 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_344 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_141 VGND VPWR sky130_fd_sc_hd__decap_12
X_5475_ _5402_/X _5406_/X _5402_/X _5406_/X _5475_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_172_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_528 VGND VPWR sky130_fd_sc_hd__decap_12
X_7214_ _7201_/X _7211_/X _7213_/Y _7214_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_4426_ _4422_/X _4424_/X _4425_/X _4426_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_67_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_678 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_509 VGND VPWR sky130_fd_sc_hd__decap_8
X_7145_ _7615_/Q _7145_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_119_1261 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_550 VGND VPWR sky130_fd_sc_hd__fill_1
X_4357_ _4830_/B _4505_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_8_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_946 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1177 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_125 VGND VPWR sky130_fd_sc_hd__decap_12
X_4288_ _4258_/X _4274_/X _4286_/X _4287_/X _4288_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_7076_ _7073_/Y _7074_/Y _7073_/Y _7074_/Y _7138_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_189_1204 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_659 VGND VPWR sky130_fd_sc_hd__decap_12
X_6027_ _6027_/A _4207_/X _6027_/C _6027_/D _6027_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_189_1248 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_512 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_865 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1240 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6929_ _7647_/Q _6929_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_2514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_559 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1126 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1186 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_261 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_581 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1156 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_373 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_970 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_384 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_928 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_631 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_472 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1074 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_166 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0_wb_clk_i clkbuf_0_wb_clk_i/X clkbuf_1_0_1_wb_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_172_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_1157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_114 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_1168 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_556 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1012 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1075 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_504 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_684 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_334 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_4483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_356 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_93 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_773 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_907 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_972 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_826 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1114 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_943 VGND VPWR sky130_fd_sc_hd__decap_3
X_5260_ _4554_/A _5123_/B _5260_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_177_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_807 VGND VPWR sky130_fd_sc_hd__decap_12
X_4211_ _4210_/X _4211_/B _4449_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_114_369 VGND VPWR sky130_fd_sc_hd__fill_2
X_5191_ _5155_/X _5159_/X _5155_/X _5159_/X _5191_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_142_689 VGND VPWR sky130_fd_sc_hd__decap_12
X_4142_ _4111_/X _4141_/X _4111_/X _4141_/X _4142_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_968 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_553 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_776 VGND VPWR sky130_fd_sc_hd__decap_12
X_4073_ _4045_/X _4046_/X _4045_/X _4046_/X _4073_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_49_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_297 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1074 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_960 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_1104 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1077 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_161 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_481 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_818 VGND VPWR sky130_fd_sc_hd__decap_12
X_7763_ _6242_/Y _5059_/A _7769_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_184_1178 VGND VPWR sky130_fd_sc_hd__decap_12
X_4975_ _4935_/X _4936_/X _4912_/X _4937_/X _4975_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_52_879 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_137 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_367 VGND VPWR sky130_fd_sc_hd__decap_12
X_6714_ _6712_/Y _6714_/B _6714_/X VGND VPWR sky130_fd_sc_hd__and2_4
XPHY_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3926_ _3926_/A _3926_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_7694_ _6675_/X _7694_/Q _7696_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_189_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_581 VGND VPWR sky130_fd_sc_hd__decap_12
X_6645_ _6636_/Y _6638_/B _6638_/X _6644_/X _6645_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_3857_ _3832_/A _3857_/B _3856_/Y _7800_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_165_737 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_428 VGND VPWR sky130_fd_sc_hd__decap_12
X_6576_ _6586_/A _6576_/B _6575_/Y _6576_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_3788_ _5128_/A _4459_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_118_642 VGND VPWR sky130_fd_sc_hd__decap_12
X_5527_ _4783_/X _4784_/X _4783_/X _4784_/X _5527_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_69_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_314 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_645 VGND VPWR sky130_fd_sc_hd__decap_8
X_5458_ _5458_/A _6006_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_117_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_656 VGND VPWR sky130_fd_sc_hd__decap_12
X_4409_ _4408_/A _4408_/B _4408_/X _4409_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_132_166 VGND VPWR sky130_fd_sc_hd__decap_12
X_5389_ _5385_/X _5388_/X _5385_/X _5388_/X _5389_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7128_ _7128_/A _7083_/X _7127_/Y _7128_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_113_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1046 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_765 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_7059_ la_data_in[86] _7060_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_59_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1056 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_813 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1237 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_548 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_98 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_152_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_654 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_520 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_52 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_721 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_715 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_202 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_940 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_409 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_910 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_984 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_697 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_678 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_964 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_452 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_306 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_986 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1096 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_713 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_724 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_938 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1077 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_139 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_843 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1104 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1115 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_818 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_643 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1001 VGND VPWR sky130_fd_sc_hd__decap_12
X_4760_ _4759_/A _4758_/X _4759_/X _4760_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XPHY_3590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_581 VGND VPWR sky130_fd_sc_hd__decap_12
X_3711_ _3711_/A _3757_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_187_873 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_682 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_715 VGND VPWR sky130_fd_sc_hd__decap_12
X_4691_ _4622_/X _4690_/X _4622_/X _4690_/X _4691_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_174_512 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_428 VGND VPWR sky130_fd_sc_hd__decap_12
X_6430_ _6412_/Y _6413_/Y _6429_/X _6431_/B VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_186_394 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_1108 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_556 VGND VPWR sky130_fd_sc_hd__decap_12
X_6361_ _6354_/A _6361_/B _6361_/C _7736_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_155_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_623 VGND VPWR sky130_fd_sc_hd__decap_8
X_5312_ _5310_/X _5311_/X _5310_/X _5311_/X _5312_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6292_ _6289_/X _6290_/Y _6291_/X _7753_/D VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_115_667 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_507 VGND VPWR sky130_fd_sc_hd__decap_12
X_5243_ _5241_/X _5242_/X _5243_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_114_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_328 VGND VPWR sky130_fd_sc_hd__decap_8
X_5174_ _5169_/X _5173_/X _5169_/X _5173_/X _5174_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_60_1005 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_1182 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_862 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1106 VGND VPWR sky130_fd_sc_hd__decap_12
X_4125_ _4122_/X _4123_/X _4131_/A _4127_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_29_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1237 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_437 VGND VPWR sky130_fd_sc_hd__decap_12
X_4056_ _4747_/B _4923_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_83_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_281 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_292 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_161 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_846 VGND VPWR sky130_fd_sc_hd__decap_8
X_7815_ _3733_/Y _7815_/Q _7810_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_307 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_306 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_654 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_318 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_879 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_329 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1095 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_507 VGND VPWR sky130_fd_sc_hd__decap_12
X_7746_ _7746_/D _7746_/Q _7746_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4958_ _4956_/X _4957_/X _4956_/X _4957_/X _4958_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_71_1134 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1262 VGND VPWR sky130_fd_sc_hd__decap_12
X_3909_ _7332_/A _3909_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_165_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1276 VGND VPWR sky130_fd_sc_hd__fill_1
X_7677_ _7677_/D _6718_/A _7658_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_177_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1118 VGND VPWR sky130_fd_sc_hd__decap_8
X_4889_ _4888_/A _4888_/B _4952_/B _4889_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_71_1189 VGND VPWR sky130_fd_sc_hd__decap_12
X_6628_ la_data_in[21] _6628_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_165_545 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_450 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_515 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_984 VGND VPWR sky130_fd_sc_hd__decap_8
X_6559_ _6595_/A _6586_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_4_739 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_634 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_291 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1074 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_678 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_65 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_912 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1252 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1274 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_562 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_1258 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_938 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_790 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_857 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1029 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_147 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_197 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_821 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_490 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_11_562 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_556 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_718 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_577 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_805 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_1253 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_98_816 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1275 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_795 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_637 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_979 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1005 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_741 VGND VPWR sky130_fd_sc_hd__decap_6
X_5930_ _5920_/Y _5921_/X _5920_/Y _5921_/X _5938_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_111_1172 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_790 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_632 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_120 VGND VPWR sky130_fd_sc_hd__fill_2
X_5861_ _5731_/A _4482_/A _5861_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_61_440 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_451 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_985 VGND VPWR sky130_fd_sc_hd__decap_12
X_7600_ _7600_/HI la_data_out[127] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_179_648 VGND VPWR sky130_fd_sc_hd__decap_12
X_4812_ _4812_/A _4814_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_107_1219 VGND VPWR sky130_fd_sc_hd__fill_1
X_5792_ _3858_/Y _4477_/A _5792_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7531_ _7531_/HI la_data_out[58] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_194_629 VGND VPWR sky130_fd_sc_hd__decap_12
X_4743_ _4743_/A _4743_/B _4743_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_203_991 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_882 VGND VPWR sky130_fd_sc_hd__decap_3
X_7462_ _7462_/HI io_out[27] VGND VPWR sky130_fd_sc_hd__conb_1
X_4674_ _4662_/X _4673_/X _4662_/X _4673_/X _4674_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_190_802 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_718 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_269 VGND VPWR sky130_fd_sc_hd__decap_3
X_6413_ la_data_in[116] _6413_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_174_364 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_887 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_910 VGND VPWR sky130_fd_sc_hd__decap_12
X_7393_ _7392_/Y _7387_/X _7773_/Q _7388_/X wbs_dat_o[27] VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1203 VGND VPWR sky130_fd_sc_hd__decap_4
X_6344_ _4126_/B _6348_/B _6347_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_179_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_740 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_954 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_208 VGND VPWR sky130_fd_sc_hd__decap_8
X_6275_ _6275_/A _6274_/X _7757_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_103_626 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_434 VGND VPWR sky130_fd_sc_hd__decap_12
X_5226_ _5212_/X _5223_/X _5224_/X _5225_/X _5226_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_97_871 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1061 VGND VPWR sky130_fd_sc_hd__decap_6
X_5157_ _5157_/A _4856_/B _5157_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_5_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_532 VGND VPWR sky130_fd_sc_hd__decap_4
X_4108_ _6095_/A _4108_/B _4211_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_99_1045 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_245 VGND VPWR sky130_fd_sc_hd__decap_12
X_5088_ _5087_/A _5087_/B _5087_/X _5088_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_84_565 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_727 VGND VPWR sky130_fd_sc_hd__decap_12
X_4039_ _4021_/X _4024_/X _4021_/X _4024_/X _4039_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_112_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_27 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_104 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_27 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_137 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_849 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_928 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_495 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_159 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1051 VGND VPWR sky130_fd_sc_hd__fill_2
X_7729_ _6448_/Y io_out[7] _7729_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_197_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1032 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_197_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1128 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_879 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_998 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_315 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_592 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_753 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_681 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_223 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1107 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1069 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_1060 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_6 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_760 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_687 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_968 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_175 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_112 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_501 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_93 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_860 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_167 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_640 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1168 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_983 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_330 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1176 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_55 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_156_364 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_875 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_868 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_280 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_740 VGND VPWR sky130_fd_sc_hd__decap_8
X_4390_ _4339_/X _4340_/X _4339_/X _4340_/X _4390_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_171_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_710 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_123 VGND VPWR sky130_fd_sc_hd__decap_12
X_6060_ _6060_/A _6060_/B _6072_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_112_445 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1220 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_871 VGND VPWR sky130_fd_sc_hd__decap_12
X_5011_ _4436_/X _4440_/X _4436_/X _4440_/X _5013_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_152_1250 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_381 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_532 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_779 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_727 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_204 VGND VPWR sky130_fd_sc_hd__decap_12
X_6962_ _7636_/Q _6962_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_19_470 VGND VPWR sky130_fd_sc_hd__fill_1
X_5913_ _5731_/A _5835_/B _5913_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_6893_ _6877_/X _6891_/X _6892_/Y _6893_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_62_760 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_985 VGND VPWR sky130_fd_sc_hd__fill_2
X_5844_ _3846_/X _5443_/B _5844_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_146_1054 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_101 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_955 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_736 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_489 VGND VPWR sky130_fd_sc_hd__decap_6
X_5775_ _5998_/A _5774_/X _5775_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_166_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_999 VGND VPWR sky130_fd_sc_hd__decap_8
X_7514_ _7514_/HI la_data_out[41] VGND VPWR sky130_fd_sc_hd__conb_1
X_4726_ _4714_/X _4724_/X _4714_/X _4724_/X _4726_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_194_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1257 VGND VPWR sky130_fd_sc_hd__decap_12
X_7445_ _7445_/HI io_out[10] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_175_684 VGND VPWR sky130_fd_sc_hd__decap_12
X_4657_ _4666_/A _4657_/B _4657_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_135_548 VGND VPWR sky130_fd_sc_hd__fill_1
X_7376_ _4794_/Y _7354_/X _7375_/X wbs_dat_o[21] VGND VPWR sky130_fd_sc_hd__o21ai_4
X_4588_ _4573_/X _4574_/X _4567_/X _4575_/X _4588_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_116_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_1033 VGND VPWR sky130_fd_sc_hd__decap_12
X_6327_ _6345_/A _6338_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_104_924 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_261 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1172 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_890 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1036 VGND VPWR sky130_fd_sc_hd__fill_1
X_6258_ _6319_/C _6249_/X _6257_/Y _6258_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_104_979 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1189 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_178 VGND VPWR sky130_fd_sc_hd__decap_12
X_5209_ _5196_/X _5206_/X _5207_/X _5208_/X _5209_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_103_489 VGND VPWR sky130_fd_sc_hd__decap_4
X_6189_ _6189_/A _6189_/B _6189_/C _6192_/A VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_40_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_705 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_362 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_215 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_259 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_719 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_944 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_112 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_443 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_977 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_145 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_426 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_758 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_138 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_353 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1122 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1193 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1245 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_905 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1199 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_803 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_814 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_863 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_727 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_226 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_708 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1273 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_387 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1246 VGND VPWR sky130_fd_sc_hd__decap_4
X_3890_ wbs_dat_i[2] _3882_/X _3891_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_32_944 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_607 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_117 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_459 VGND VPWR sky130_fd_sc_hd__decap_8
X_5560_ _5552_/X _5553_/X _5558_/X _5559_/X _5560_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_129_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_4511_ _4503_/X _4507_/X _4503_/X _4507_/X _4511_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_106_1093 VGND VPWR sky130_fd_sc_hd__decap_12
X_5491_ _5489_/X _5490_/X _5491_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_117_548 VGND VPWR sky130_fd_sc_hd__fill_1
X_7230_ _7193_/X _7228_/X _7229_/Y _7230_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_7_182 VGND VPWR sky130_fd_sc_hd__fill_1
X_4442_ _4386_/X _4441_/X _4443_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_172_654 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_879 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_172_676 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_900 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_518 VGND VPWR sky130_fd_sc_hd__fill_1
X_7161_ la_data_in[104] _7161_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_144_389 VGND VPWR sky130_fd_sc_hd__decap_8
X_4373_ _4368_/X _4372_/B _4372_/X _4373_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_98_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1206 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_592 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_955 VGND VPWR sky130_fd_sc_hd__fill_2
X_6112_ _4210_/B _6112_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_99_966 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_540 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_977 VGND VPWR sky130_fd_sc_hd__decap_12
X_7092_ _7043_/Y _7044_/Y _7045_/X _7091_/X _7092_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_59_819 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_307 VGND VPWR sky130_fd_sc_hd__decap_12
X_6043_ wb_rst_i _6044_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_67_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_448 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1008 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_1121 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1199 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1143 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_321 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1116 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6945_ la_data_in[72] _6945_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_3419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_782 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_410 VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_2_2_0_wb_clk_i clkbuf_1_1_1_wb_clk_i/X clkbuf_2_2_1_wb_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_6876_ _6833_/A _6832_/Y _6833_/X _6875_/X _6876_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XPHY_2729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_938 VGND VPWR sky130_fd_sc_hd__decap_8
X_5827_ _3901_/X _4295_/Y _5827_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_23_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_605 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1081 VGND VPWR sky130_fd_sc_hd__decap_8
X_5758_ _5747_/X _5748_/X _5747_/X _5748_/X _5758_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_124_1171 VGND VPWR sky130_fd_sc_hd__decap_12
X_4709_ _4692_/X _4706_/X _4707_/X _4708_/X _4709_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_185_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_5689_ _5687_/X _5688_/X _5689_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_108_548 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1117 VGND VPWR sky130_fd_sc_hd__decap_12
X_7428_ io_oeb[23] _7428_/LO VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_159_1245 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_698 VGND VPWR sky130_fd_sc_hd__decap_4
X_7359_ _5277_/Y _7355_/X _7358_/X wbs_dat_o[16] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_116_581 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_798 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_971 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_513 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_855 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_74 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_708 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_96 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_4654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_527 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_922 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_398 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_916 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_999 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_436 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_498 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1252 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_662 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_418 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_963 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_631 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_440 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_653 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_551 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_616 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_150_882 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_413 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_947 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1250 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_611 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_768 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_811 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_833 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1030 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_568 VGND VPWR sky130_fd_sc_hd__decap_12
X_4991_ _4990_/X _4991_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_6730_ _7673_/Q _6730_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_51_538 VGND VPWR sky130_fd_sc_hd__decap_8
X_3942_ _4959_/A _4078_/B _3942_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_189_562 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_724 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1065 VGND VPWR sky130_fd_sc_hd__decap_3
X_6661_ _6602_/X _6667_/B _6661_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_3873_ wbs_dat_i[4] _3848_/B _3874_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_189_595 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1046 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_1166 VGND VPWR sky130_fd_sc_hd__decap_12
X_5612_ _5605_/X _5611_/X _5605_/X _5611_/X _5612_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_104_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_273 VGND VPWR sky130_fd_sc_hd__decap_12
X_6592_ _7700_/Q la_data_in[2] _6530_/X _6592_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_192_727 VGND VPWR sky130_fd_sc_hd__decap_12
X_5543_ _5537_/X _5538_/X _5536_/X _5539_/X _5543_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_145_632 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_857 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_480 VGND VPWR sky130_fd_sc_hd__decap_4
X_5474_ _5472_/X _5473_/X _5474_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_117_356 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_367 VGND VPWR sky130_fd_sc_hd__decap_12
X_7213_ _7201_/X _7211_/X _7212_/X _7213_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_145_698 VGND VPWR sky130_fd_sc_hd__decap_12
X_4425_ _4422_/X _4424_/X _4425_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_172_495 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_1172 VGND VPWR sky130_fd_sc_hd__decap_8
X_7144_ _7142_/Y _7143_/Y _7142_/Y _7143_/Y _7144_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_63_1014 VGND VPWR sky130_fd_sc_hd__decap_12
X_4356_ _4820_/A _4498_/B _4359_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_87_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_871 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1273 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_936 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1006 VGND VPWR sky130_fd_sc_hd__fill_1
X_7075_ _7618_/Q la_data_in[80] _7077_/A VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_87_958 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1189 VGND VPWR sky130_fd_sc_hd__fill_1
X_4287_ _4258_/X _4274_/X _4258_/X _4274_/X _4287_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_101_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_137 VGND VPWR sky130_fd_sc_hd__decap_12
X_6026_ _4449_/A _6025_/X _6027_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_39_351 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_524 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_855 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_708 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_398 VGND VPWR sky130_fd_sc_hd__decap_6
X_6928_ _6926_/Y _6927_/Y _6926_/Y _6927_/Y _6993_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_2515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_56 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_831 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_27 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_914 VGND VPWR sky130_fd_sc_hd__fill_1
X_6859_ la_data_in[49] _6859_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_1825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_273 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_593 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_424 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_621 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_98 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_440 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_782 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_601 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_484 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_612 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1231 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_551 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_155 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_800 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_811 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_663 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_365 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1087 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_516 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_368 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_200 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_785 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_582 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_886 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_727 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_429 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_790 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_1093 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_760 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_451 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_911 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_984 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_838 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1126 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_337 VGND VPWR sky130_fd_sc_hd__fill_1
X_4210_ _4208_/X _4210_/B _4210_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_130_819 VGND VPWR sky130_fd_sc_hd__decap_4
X_5190_ _5185_/X _5189_/X _5188_/X _5190_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_69_936 VGND VPWR sky130_fd_sc_hd__fill_1
X_4141_ _4112_/X _4129_/X _4130_/X _4140_/X _4141_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_110_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_755 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_232 VGND VPWR sky130_fd_sc_hd__decap_12
X_4072_ _4048_/X _4060_/X _4048_/X _4060_/X _4072_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_565 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_788 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_107 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1233 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_1067 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1116 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_825 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_696 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_173 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_387 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_184 VGND VPWR sky130_fd_sc_hd__decap_8
X_4974_ _4962_/X _4973_/X _4962_/X _4973_/X _4974_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7762_ _7762_/D _7762_/Q _7769_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_3925_ _3689_/A _3928_/A _3926_/A VGND VPWR sky130_fd_sc_hd__and2_4
X_6713_ la_data_in[45] _6714_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_51_379 VGND VPWR sky130_fd_sc_hd__decap_12
X_7693_ _6678_/X _6609_/A _7696_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_211_149 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_245 VGND VPWR sky130_fd_sc_hd__decap_4
X_6644_ _6639_/Y _6640_/Y _6643_/X _6644_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_32_593 VGND VPWR sky130_fd_sc_hd__decap_12
X_3856_ wbs_dat_i[6] _3848_/B _3856_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_165_716 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_407 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_587 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_6575_ _6575_/A _6546_/X _6575_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_3787_ _4553_/A _5128_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_5526_ _5315_/X _5316_/X _5314_/X _5317_/X _5526_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_145_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_900 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_1245 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1215 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_410 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_849 VGND VPWR sky130_fd_sc_hd__decap_12
X_5457_ _5455_/X _6006_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_59_28 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_668 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_808 VGND VPWR sky130_fd_sc_hd__decap_12
X_4408_ _4408_/A _4408_/B _4408_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_133_679 VGND VPWR sky130_fd_sc_hd__decap_8
X_5388_ _5386_/X _5387_/X _5386_/X _5387_/X _5388_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_87_700 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_178 VGND VPWR sky130_fd_sc_hd__decap_12
X_7127_ _7083_/A _7083_/B _7127_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_87_733 VGND VPWR sky130_fd_sc_hd__decap_12
X_4339_ _4337_/X _4338_/X _4337_/X _4338_/X _4339_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_87_777 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1069 VGND VPWR sky130_fd_sc_hd__decap_12
X_7058_ _7058_/A _7058_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_189_1013 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_276 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_1191 VGND VPWR sky130_fd_sc_hd__decap_12
X_6009_ _5334_/B _6005_/Y _6008_/Y _6010_/B VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_101_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_354 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_123 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_471 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1249 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1219 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_335 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_346 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_666 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1090 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_64 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_891 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_733 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_502 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_683 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_587 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_418 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_269 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_996 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1020 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_998 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1023 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_83 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1089 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_674 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1127 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1191 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_655 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_379 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1013 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_841 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3710_ _3710_/A _6323_/A _3711_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_159_554 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1163 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1166 VGND VPWR sky130_fd_sc_hd__decap_12
X_4690_ _4675_/X _4689_/X _4675_/X _4689_/X _4690_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_41_390 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_727 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_568 VGND VPWR sky130_fd_sc_hd__decap_12
X_6360_ wbs_dat_i[6] _6349_/B _6361_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_127_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_3 VGND VPWR sky130_fd_sc_hd__decap_4
X_5311_ _5160_/X _5166_/X _5154_/X _5167_/X _5311_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_142_410 VGND VPWR sky130_fd_sc_hd__decap_12
X_6291_ _5845_/Y _6256_/B _3743_/A _6291_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_143_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_808 VGND VPWR sky130_fd_sc_hd__decap_12
X_5242_ _4716_/A _4460_/B _5242_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_130_616 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1142 VGND VPWR sky130_fd_sc_hd__fill_1
X_5173_ _5172_/A _5172_/B _5172_/X _5173_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_4124_ _4122_/X _4123_/X _4131_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_84_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1028 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_874 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1118 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1249 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1080 VGND VPWR sky130_fd_sc_hd__decap_12
X_4055_ _4624_/B _4747_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_56_449 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_260 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_685 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_173 VGND VPWR sky130_fd_sc_hd__fill_1
X_7814_ _3741_/Y _7814_/Q _7810_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_51_121 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_308 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_319 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_666 VGND VPWR sky130_fd_sc_hd__decap_8
X_4957_ _4905_/X _4906_/X _4904_/X _4957_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_7745_ _6329_/Y _3919_/A _7810_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_75_1271 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1252 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_1146 VGND VPWR sky130_fd_sc_hd__decap_12
X_3908_ _7338_/A _6042_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_4888_ _4888_/A _4888_/B _4952_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7676_ _7676_/D _7676_/Q _7707_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_162_1274 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_165_513 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_727 VGND VPWR sky130_fd_sc_hd__decap_6
X_3839_ _3759_/A _3848_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_6627_ _6627_/A _6627_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_193_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_952 VGND VPWR sky130_fd_sc_hd__decap_12
X_6558_ _6885_/A _6556_/Y _6558_/C _6558_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_69_1031 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_398 VGND VPWR sky130_fd_sc_hd__decap_12
X_5509_ _5506_/X _5508_/X _5506_/X _5508_/X _5509_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_180_549 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_6489_ _7714_/Q la_data_in[112] _6489_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_105_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_44 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_77 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_627 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_1029 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1242 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_906 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_928 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_265 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_585 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1275 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_611 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_121 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1019 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_806 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_959 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_74 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_154 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1002 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1024 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_51 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_62 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_585 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_73 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1030 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1090 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_589 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1101 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_292 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1145 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1148 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_649 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_563 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1017 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_449 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1181 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_685 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_931 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1203 VGND VPWR sky130_fd_sc_hd__decap_12
X_5860_ _3875_/Y _4477_/A _5860_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_206_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_655 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1116 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_80 VGND VPWR sky130_fd_sc_hd__decap_12
X_4811_ _4603_/X _4620_/X _4588_/X _4621_/X _4811_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_61_463 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_907 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_997 VGND VPWR sky130_fd_sc_hd__decap_8
X_5791_ _5786_/X _5790_/X _5789_/X _5791_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_34_699 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_891 VGND VPWR sky130_fd_sc_hd__decap_3
X_4742_ _4742_/A _3930_/A _4742_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7530_ _7530_/HI la_data_out[57] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_14_390 VGND VPWR sky130_fd_sc_hd__decap_6
X_7461_ _7461_/HI io_out[26] VGND VPWR sky130_fd_sc_hd__conb_1
X_4673_ _4663_/X _4670_/X _4671_/X _4672_/X _4673_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_175_855 VGND VPWR sky130_fd_sc_hd__decap_12
X_6412_ _6412_/A _6412_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_190_814 VGND VPWR sky130_fd_sc_hd__decap_8
X_7392_ io_in[33] _7392_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_174_376 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_922 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_398 VGND VPWR sky130_fd_sc_hd__decap_12
X_6343_ _6350_/A _6343_/B _6342_/Y _6343_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_127_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_966 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1226 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_763 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_605 VGND VPWR sky130_fd_sc_hd__decap_4
X_6274_ _5639_/Y _6091_/X _6208_/A _6274_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_89_828 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_638 VGND VPWR sky130_fd_sc_hd__decap_3
X_5225_ _5212_/X _5223_/X _5212_/X _5223_/X _5225_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_170_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1131 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_850 VGND VPWR sky130_fd_sc_hd__decap_4
X_5156_ _5171_/A _4854_/B _5156_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_69_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_213 VGND VPWR sky130_fd_sc_hd__fill_1
X_4107_ _4102_/A _4206_/A _4102_/A _4206_/A _4108_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_5087_ _5087_/A _5087_/B _5087_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_56_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_577 VGND VPWR sky130_fd_sc_hd__decap_3
X_4038_ _7783_/Q _4038_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_38_983 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_739 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_121 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_964 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_105 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_761 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_806 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_116 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_154 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_127 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VPWR sky130_fd_sc_hd__decap_3
X_5989_ _5883_/X _6280_/A _5988_/X _5990_/B VGND VPWR sky130_fd_sc_hd__o21a_4
XPHY_149 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_619 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_349 VGND VPWR sky130_fd_sc_hd__decap_12
X_7728_ _7728_/D _7728_/Q _7785_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_138_513 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1093 VGND VPWR sky130_fd_sc_hd__fill_2
X_7659_ _6901_/X _6834_/A _7658_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_197_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_292 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_465 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_796 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_582 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_765 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_776 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_693 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_1026 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_235 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1119 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_471 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_611 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_227 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_547 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_482 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_633 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_7 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_772 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_699 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_468 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_647 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_124 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1114 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_991 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_524 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_872 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_179 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_894 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_23 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1106 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_708 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_995 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_376 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_549 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_292 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_379 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_4_0_wb_clk_i clkbuf_2_2_1_wb_clk_i/X clkbuf_4_9_0_wb_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_194_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_880 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1062 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_722 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_457 VGND VPWR sky130_fd_sc_hd__fill_1
X_5010_ _4992_/X _5008_/X _5005_/X _5009_/X _5012_/A VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_140_788 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_883 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_511 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_393 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_758 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_555 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_886 VGND VPWR sky130_fd_sc_hd__decap_12
X_6961_ _6959_/Y _6960_/Y _6961_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_81_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_739 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_216 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1094 VGND VPWR sky130_fd_sc_hd__decap_12
X_5912_ _5894_/Y _5895_/X _5894_/Y _5895_/X _5912_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6892_ _6877_/X _6891_/X _6811_/X _6892_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_5843_ _5833_/X _5836_/X _5843_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_195_906 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_1066 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_113 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_928 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_135 VGND VPWR sky130_fd_sc_hd__decap_12
X_5774_ _5767_/X _5772_/X _5774_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_188_980 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1252 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_166_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_7513_ _7513_/HI la_data_out[40] VGND VPWR sky130_fd_sc_hd__conb_1
X_4725_ _4472_/X _4473_/X _4472_/X _4473_/X _4725_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_147_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1269 VGND VPWR sky130_fd_sc_hd__decap_8
X_4656_ _4656_/A _4666_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_7444_ _7444_/HI io_out[9] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_148_899 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_335 VGND VPWR sky130_fd_sc_hd__fill_1
X_4587_ _4545_/X _4586_/X _4545_/X _4586_/X _4587_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7375_ _4793_/A _7370_/X _7374_/Y _7364_/X _7375_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_6326_ _6340_/A _6345_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_1_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_699 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_1045 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_733 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_947 VGND VPWR sky130_fd_sc_hd__decap_12
X_6257_ _5779_/X _6248_/X _6257_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_67_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_5208_ _5196_/X _5206_/X _5196_/X _5206_/X _5208_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_131_788 VGND VPWR sky130_fd_sc_hd__decap_4
X_6188_ _4884_/X _6186_/Y _6189_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_130_276 VGND VPWR sky130_fd_sc_hd__decap_12
X_5139_ _5157_/A _4854_/B _5140_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_85_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_886 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_897 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_65 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1275 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_956 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_124 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_365 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_505 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_685 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1172 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_879 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_180_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_880 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_699 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_722 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_1265 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_593 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_917 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_265 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_831 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_826 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_875 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_83 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1201 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_739 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_216 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_845 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_238 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1234 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_558 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_964 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_733 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_761 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_744 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1127 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1209 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_129 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1080 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1001 VGND VPWR sky130_fd_sc_hd__decap_4
X_4510_ _4496_/X _4509_/X _4496_/X _4509_/X _4510_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_129_354 VGND VPWR sky130_fd_sc_hd__decap_12
X_5490_ _3813_/X _4782_/B _5490_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1004 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_171_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_633 VGND VPWR sky130_fd_sc_hd__decap_8
X_4441_ _4387_/X _4439_/X _4436_/X _4440_/X _4441_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_176_1037 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_912 VGND VPWR sky130_fd_sc_hd__decap_3
X_7160_ _7160_/A _7160_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_172_688 VGND VPWR sky130_fd_sc_hd__decap_12
X_4372_ _4368_/X _4372_/B _4372_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_153_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_422 VGND VPWR sky130_fd_sc_hd__decap_12
X_6111_ _6185_/A _6111_/B _7784_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_113_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1218 VGND VPWR sky130_fd_sc_hd__fill_2
X_7091_ _7048_/A _7048_/B _7048_/X _7090_/X _7091_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_101_906 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_552 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_989 VGND VPWR sky130_fd_sc_hd__decap_6
X_6042_ _6042_/A _3909_/Y _3910_/Y _6058_/B _6050_/B VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_101_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_319 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1040 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1155 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_508 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_1166 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_333 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1128 VGND VPWR sky130_fd_sc_hd__fill_1
X_6944_ _7642_/Q _6944_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_19_290 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_912 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6875_ _6834_/Y _6835_/Y _6874_/X _6875_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_179_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_794 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_714 VGND VPWR sky130_fd_sc_hd__decap_12
X_5826_ _5786_/X _5790_/X _5786_/X _5790_/X _5826_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_210_523 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_989 VGND VPWR sky130_fd_sc_hd__decap_12
X_5757_ _5753_/X _5756_/X _5753_/X _5756_/X _5757_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_120_1014 VGND VPWR sky130_fd_sc_hd__decap_12
X_4708_ _4692_/X _4706_/X _4692_/X _4706_/X _4708_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_163_600 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_825 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_1183 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_611 VGND VPWR sky130_fd_sc_hd__fill_1
X_5688_ _3843_/A _4820_/B _5688_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_147_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1099 VGND VPWR sky130_fd_sc_hd__decap_8
X_7427_ io_oeb[22] _7427_/LO VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_120_1069 VGND VPWR sky130_fd_sc_hd__decap_4
X_4639_ _5128_/A _4624_/B _4639_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_190_441 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_964 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_997 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1093 VGND VPWR sky130_fd_sc_hd__decap_12
X_7358_ _3773_/X _7349_/X _7356_/Y _7387_/A _7358_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_104_711 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_6309_ _5974_/A _5973_/X _5974_/A _5973_/X _6309_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_104_755 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_232 VGND VPWR sky130_fd_sc_hd__decap_12
X_7289_ _5176_/A _7262_/X _7288_/X _7289_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_131_574 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_820 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1004 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_609 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1143 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_983 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_300 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_694 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_306 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_32 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_867 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1050 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_934 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_501 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_928 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_641 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1250 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_1182 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_296 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_920 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_357 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_665 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1032 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_563 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_601 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_875 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_672 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_620 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_845 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_141 VGND VPWR sky130_fd_sc_hd__decap_12
X_4990_ _4983_/X _4989_/X _4990_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_205_851 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_1011 VGND VPWR sky130_fd_sc_hd__decap_8
X_3941_ _4164_/B _4078_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_56_1022 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_794 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1097 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_3872_ _5176_/A _3838_/B _3874_/B VGND VPWR sky130_fd_sc_hd__and2_4
X_6660_ _6605_/A _6605_/B _6605_/X _6659_/X _6667_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_176_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_263 VGND VPWR sky130_fd_sc_hd__fill_1
X_5611_ _5606_/X _5610_/X _5609_/X _5611_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_108_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_950 VGND VPWR sky130_fd_sc_hd__decap_12
X_6591_ _6537_/X _6589_/X _6590_/Y _6591_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_5542_ _5522_/X _5531_/X _5540_/X _5541_/X _5542_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_192_739 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_825 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_993 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_493 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_184 VGND VPWR sky130_fd_sc_hd__decap_12
X_5473_ _5216_/A _4747_/B _5473_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_118_869 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_154 VGND VPWR sky130_fd_sc_hd__decap_12
X_4424_ _4561_/A _4903_/B _4424_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7212_ _6068_/A _7212_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_117_379 VGND VPWR sky130_fd_sc_hd__decap_12
X_4355_ _4613_/B _4498_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_7143_ la_data_in[110] _7143_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_113_541 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_775 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1026 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_563 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_883 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_263 VGND VPWR sky130_fd_sc_hd__decap_12
X_7074_ la_data_in[81] _7074_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_58_105 VGND VPWR sky130_fd_sc_hd__decap_6
X_4286_ _4282_/X _4285_/X _4282_/X _4285_/X _4286_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_100_202 VGND VPWR sky130_fd_sc_hd__decap_12
X_6025_ _4450_/X _4451_/X _6025_/C _6024_/Y _6025_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_101_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_149 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_363 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_536 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_642 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_889 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_506 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6927_ la_data_in[78] _6927_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_3239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_731 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_703 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_68 VGND VPWR sky130_fd_sc_hd__decap_12
X_6858_ _7651_/Q _6858_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_1815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5809_ _5805_/X _5806_/X _5807_/Y _5808_/X _5809_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XPHY_1848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_948 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6789_ _6765_/X _6788_/X _6785_/X _6789_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_167_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_566 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_436 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1010 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_699 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_794 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_891 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_1240 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_635 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_861 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_145 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1243 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_563 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_679 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_883 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_178 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_469 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_981 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_791 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_141 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_528 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_51 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1069 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_550 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_285 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_245 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_739 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_666 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_923 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_996 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_1059 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1018 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1149 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_701 VGND VPWR sky130_fd_sc_hd__fill_1
X_4140_ _4132_/X _4139_/X _4140_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_150_691 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_544 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_907 VGND VPWR sky130_fd_sc_hd__decap_8
X_4071_ _4062_/X _4063_/X _4062_/X _4063_/X _4092_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_84_918 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_609 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_431 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_577 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_428 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_620 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1250 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1212 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_141 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1128 VGND VPWR sky130_fd_sc_hd__fill_1
X_7761_ _7761_/D _5383_/A _7758_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4973_ _4971_/X _4972_/X _4971_/X _4972_/X _4973_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_211_106 VGND VPWR sky130_fd_sc_hd__decap_12
X_6712_ _7679_/Q _6712_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_3924_ _3949_/B _3924_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_7692_ _6681_/X _6612_/A _7696_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_6643_ _6705_/A _6642_/X _6643_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_3855_ _5137_/A _3838_/B _3857_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_165_728 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_419 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_599 VGND VPWR sky130_fd_sc_hd__decap_8
X_3786_ _3786_/A _4553_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_6574_ _6548_/X _6571_/X _6573_/Y _6574_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_164_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_110 VGND VPWR sky130_fd_sc_hd__decap_12
X_5525_ _5307_/X _5308_/X _5306_/X _5309_/X _5525_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_195_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_912 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_794 VGND VPWR sky130_fd_sc_hd__decap_12
X_5456_ _5392_/X _5393_/X _5392_/X _5393_/X _5458_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_4407_ _4847_/A _4461_/B _4408_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_161_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_550 VGND VPWR sky130_fd_sc_hd__decap_4
X_5387_ _5277_/Y _5278_/X _5277_/Y _5278_/X _5387_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_87_712 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_403 VGND VPWR sky130_fd_sc_hd__decap_12
X_7126_ _7084_/X _7124_/X _7125_/Y _7624_/D VGND VPWR sky130_fd_sc_hd__o21a_4
X_4338_ _5304_/A _4546_/B _4338_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_87_745 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_190 VGND VPWR sky130_fd_sc_hd__decap_12
X_4269_ _4269_/A _4268_/X _4269_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7057_ _7057_/A _7057_/B _7057_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_87_789 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_1025 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_6008_ _6008_/A _6008_/B _6008_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_28_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_300 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_141 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_483 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_27 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1050 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_3058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_500 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_358 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_678 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_509 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_32 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1031 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_544 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_76 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_745 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_886 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_705 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_514 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_695 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1250 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_611 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_215 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_558 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_1245 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_288 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_761 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_772 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_614 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_809 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_977 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1051 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_487 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_498 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1035 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_95 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_36 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_47 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_50 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_344 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_623 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_837 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_1139 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_196 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_667 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_4293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1172 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_1142 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_1025 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_190 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1175 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_208 VGND VPWR sky130_fd_sc_hd__decap_12
X_5310_ _5306_/X _5309_/X _5306_/X _5309_/X _5310_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6290_ _5984_/Y _6288_/X _6101_/X _6290_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_155_794 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_934 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_422 VGND VPWR sky130_fd_sc_hd__decap_12
X_5241_ _4741_/A _4461_/B _5241_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_170_764 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_143_989 VGND VPWR sky130_fd_sc_hd__decap_12
X_5172_ _5172_/A _5172_/B _5172_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_96_520 VGND VPWR sky130_fd_sc_hd__decap_6
X_4123_ _3738_/X _4123_/B _4123_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_64_1187 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_907 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_288 VGND VPWR sky130_fd_sc_hd__decap_12
X_4054_ _4054_/A _4624_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_110_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1092 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_272 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_910 VGND VPWR sky130_fd_sc_hd__decap_12
X_7813_ _3751_/Y _7813_/Q _7810_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_483 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_697 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_309 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_7744_ _7744_/D _3928_/A _7810_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4956_ _4426_/X _4428_/X _4426_/X _4428_/X _4956_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_101_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_998 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_853 VGND VPWR sky130_fd_sc_hd__fill_1
X_3907_ _3866_/X _3907_/B _3907_/C _7794_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_20_520 VGND VPWR sky130_fd_sc_hd__decap_12
X_7675_ _6793_/X _7675_/Q _7756_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4887_ _4887_/A _4825_/X _4888_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_178_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_300 VGND VPWR sky130_fd_sc_hd__decap_12
X_6626_ _6624_/Y _6625_/Y _6626_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_3838_ _5420_/A _3838_/B _3841_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_193_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_249 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_964 VGND VPWR sky130_fd_sc_hd__decap_12
X_6557_ la_data_in[15] _6556_/B _6558_/C VGND VPWR sky130_fd_sc_hd__and2_4
X_3769_ _3769_/A _3767_/X _3768_/Y _3769_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_5508_ _5507_/A _5445_/Y _5507_/X _5508_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_134_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_23 VGND VPWR sky130_fd_sc_hd__decap_8
X_6488_ _6466_/X _6488_/B _6487_/Y _6488_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_105_135 VGND VPWR sky130_fd_sc_hd__decap_12
X_5439_ _5401_/X _5418_/X _5401_/X _5418_/X _5439_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_117_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_89 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_7109_ _7092_/X _7107_/X _7108_/Y _7630_/D VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_101_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_597 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_770 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_461 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_837 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_6_0_wb_clk_i clkbuf_4_7_0_wb_clk_i/A _7758_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_188_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_133 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_86 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_853 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1036 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_171 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_227 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_85 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_597 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_441 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1132 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_485 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1097 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_422 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_1113 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1067 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_764 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_306 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_959 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_691 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_661 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_501 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_575 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1002 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1103 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_697 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_943 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_667 VGND VPWR sky130_fd_sc_hd__decap_12
X_4810_ _4581_/X _4583_/X _4580_/Y _4584_/X _4810_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XPHY_4090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5790_ _5789_/A _5789_/B _5789_/X _5790_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_21_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_919 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_330 VGND VPWR sky130_fd_sc_hd__decap_12
X_4741_ _4741_/A _4665_/B _4741_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_187_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_300 VGND VPWR sky130_fd_sc_hd__decap_12
X_7460_ _7460_/HI io_out[25] VGND VPWR sky130_fd_sc_hd__conb_1
X_4672_ _4663_/X _4670_/X _4663_/X _4670_/X _4672_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_174_322 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_867 VGND VPWR sky130_fd_sc_hd__decap_12
X_6411_ _6409_/Y _6410_/Y _6409_/Y _6410_/Y _6431_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_31_1131 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_1035 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_1191 VGND VPWR sky130_fd_sc_hd__decap_12
X_7391_ _7390_/Y _7387_/X _4886_/A _7388_/X wbs_dat_o[26] VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_190_837 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_388 VGND VPWR sky130_fd_sc_hd__decap_8
X_6342_ wbs_dat_i[11] _6338_/B _6342_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_116_934 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_411 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_807 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_978 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1238 VGND VPWR sky130_fd_sc_hd__decap_12
X_6273_ _6240_/A _6273_/B _6273_/C _6275_/A VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_143_775 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_306 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_5224_ _5116_/X _5117_/X _5116_/X _5117_/X _5224_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_142_296 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_1143 VGND VPWR sky130_fd_sc_hd__decap_12
X_5155_ _4695_/A _4852_/B _5155_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_111_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_428 VGND VPWR sky130_fd_sc_hd__decap_12
X_4106_ _3996_/X _4031_/X _4032_/X _4206_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
X_5086_ _4749_/A _4596_/B _5087_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_99_1036 VGND VPWR sky130_fd_sc_hd__fill_1
X_4037_ _4032_/X _4034_/B _4036_/Y _6028_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_56_269 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_770 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_995 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1209 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_106 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_818 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_128 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_198_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_166 VGND VPWR sky130_fd_sc_hd__decap_12
X_5988_ _5858_/X _5988_/B _5988_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_139 VGND VPWR sky130_fd_sc_hd__decap_3
X_7727_ _6453_/X _7727_/Q _7785_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4939_ _4871_/X _4872_/X _4838_/X _4873_/X _4939_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_166_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_834 VGND VPWR sky130_fd_sc_hd__decap_12
X_7658_ _6903_/X _6837_/A _7658_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_177_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1056 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_11 VGND VPWR sky130_fd_sc_hd__fill_2
X_6609_ _6609_/A _6611_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_197_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_901 VGND VPWR sky130_fd_sc_hd__decap_12
X_7589_ _7589_/HI la_data_out[116] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_181_826 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1108 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_794 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_1160 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_1171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1005 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_41 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_494 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_740 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_8 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_784 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1142 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_136 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_840 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_672 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1126 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_884 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_867 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1118 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_889 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_506 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_388 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_775 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1074 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_948 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_734 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1135 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_810 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_361 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_567 VGND VPWR sky130_fd_sc_hd__decap_12
X_6960_ la_data_in[67] _6960_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_94_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_228 VGND VPWR sky130_fd_sc_hd__decap_12
X_5911_ _5886_/X _5904_/X _5905_/X _5911_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_207_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_943 VGND VPWR sky130_fd_sc_hd__decap_8
X_6891_ _6825_/A la_data_in[60] _6827_/X _6891_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_62_740 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_425 VGND VPWR sky130_fd_sc_hd__fill_2
X_5842_ _5783_/X _5802_/X _5803_/X _5842_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_22_626 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1029 VGND VPWR sky130_fd_sc_hd__decap_8
X_5773_ _5767_/X _5772_/X _5998_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_21_147 VGND VPWR sky130_fd_sc_hd__decap_12
X_7512_ _7512_/HI la_data_out[39] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_188_992 VGND VPWR sky130_fd_sc_hd__decap_12
X_4724_ _4715_/X _4721_/X _4722_/X _4723_/X _4724_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_159_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_480 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_681 VGND VPWR sky130_fd_sc_hd__decap_12
X_7443_ _7443_/HI io_out[8] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_174_141 VGND VPWR sky130_fd_sc_hd__decap_12
X_4655_ _4655_/A _4666_/B _4655_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_107_208 VGND VPWR sky130_fd_sc_hd__decap_12
X_7374_ io_in[27] _7374_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_200_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_731 VGND VPWR sky130_fd_sc_hd__decap_8
X_4586_ _4579_/X _4585_/X _4579_/X _4585_/X _4586_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_116_742 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_667 VGND VPWR sky130_fd_sc_hd__decap_12
X_6325_ _3924_/X _6334_/B _6329_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_143_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_519 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1057 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1019 VGND VPWR sky130_fd_sc_hd__decap_12
X_6256_ _5507_/A _6256_/B _6256_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_104_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_756 VGND VPWR sky130_fd_sc_hd__decap_8
X_5207_ _5149_/X _5150_/X _5149_/X _5150_/X _5207_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6187_ _4884_/X _6186_/Y _6189_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_57_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_692 VGND VPWR sky130_fd_sc_hd__decap_12
X_5138_ _4718_/A _4856_/B _5140_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_111_480 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_269 VGND VPWR sky130_fd_sc_hd__decap_12
X_5069_ _5069_/A _5294_/B _5069_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_45_729 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_910 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_83_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_943 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_751 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_44 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_604 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_77 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_581 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_497 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_968 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_166_697 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_1230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1067 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_607 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_929 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_95 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_898 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_375 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1213 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1246 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1253 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_924 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_784 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_756 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_581 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_907 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_456 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_288 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_480 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_489 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_1092 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_631 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_670 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_1013 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_141 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_483 VGND VPWR sky130_fd_sc_hd__decap_12
X_4440_ _4387_/X _4439_/X _4387_/X _4439_/X _4440_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_7_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1049 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_550 VGND VPWR sky130_fd_sc_hd__decap_12
X_4371_ _4369_/X _4370_/X _4369_/X _4370_/X _4372_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_208_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_935 VGND VPWR sky130_fd_sc_hd__decap_12
X_6110_ _6106_/X _6107_/X _6108_/X _7784_/Q _6109_/X _6111_/B VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_98_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_520 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_434 VGND VPWR sky130_fd_sc_hd__decap_12
X_7090_ _7049_/Y _7050_/Y _7118_/B _7090_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_113_745 VGND VPWR sky130_fd_sc_hd__decap_12
X_6041_ _6029_/X _6034_/X _6139_/A _6058_/B VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_140_564 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1090 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1074 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_364 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_239 VGND VPWR sky130_fd_sc_hd__decap_8
X_6943_ _6941_/Y _6942_/Y _6941_/Y _6942_/Y _7008_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_208_882 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_367 VGND VPWR sky130_fd_sc_hd__decap_12
X_6874_ _6874_/A _6873_/X _6874_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_2709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_721 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_581 VGND VPWR sky130_fd_sc_hd__decap_12
X_5825_ _5798_/X _5799_/X _5798_/X _5799_/X _5825_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_23_968 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_726 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_167_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_535 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_467 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_618 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_1181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_478 VGND VPWR sky130_fd_sc_hd__decap_12
X_5756_ _5745_/X _5755_/X _5745_/X _5755_/X _5756_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_148_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_579 VGND VPWR sky130_fd_sc_hd__fill_1
X_4707_ _4577_/X _4578_/X _4577_/X _4578_/X _4707_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_176_984 VGND VPWR sky130_fd_sc_hd__decap_12
X_5687_ _4680_/A _5301_/B _5687_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_120_1026 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1037 VGND VPWR sky130_fd_sc_hd__decap_12
X_7426_ io_oeb[21] _7426_/LO VGND VPWR sky130_fd_sc_hd__conb_1
X_4638_ _4623_/X _4637_/X _4623_/X _4637_/X _4638_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_147_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_190_453 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_818 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_509 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_1149 VGND VPWR sky130_fd_sc_hd__decap_8
X_7357_ _7265_/X _7387_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_162_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_68 VGND VPWR sky130_fd_sc_hd__decap_12
X_4569_ _4519_/A _4569_/B _4569_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_2_828 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_839 VGND VPWR sky130_fd_sc_hd__decap_8
X_6308_ _5946_/A _6308_/B _6308_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_7288_ _7288_/A _7300_/B _7288_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_6239_ _6198_/A _6238_/B _6240_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_89_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1155 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_995 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1248 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_537 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_1259 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_44 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_879 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_773 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_784 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_581 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1084 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_416 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_1005 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_653 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_303 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_932 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_678 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1052 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_520 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_1082 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_862 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_715 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_575 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_726 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_624 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_632 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1050 VGND VPWR sky130_fd_sc_hd__decap_12
X_3940_ _4328_/B _4164_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_16_250 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1020 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_890 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_732 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_220 VGND VPWR sky130_fd_sc_hd__decap_12
X_3871_ _5348_/A _5176_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_147_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_428 VGND VPWR sky130_fd_sc_hd__decap_12
X_5610_ _5607_/X _5608_/X _5609_/X _5610_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_6590_ _6537_/X _6589_/X _6572_/X _6590_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_83_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_962 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_297 VGND VPWR sky130_fd_sc_hd__decap_8
X_5541_ _5522_/X _5531_/X _5522_/X _5531_/X _5541_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_118_815 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_984 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_770 VGND VPWR sky130_fd_sc_hd__fill_1
X_5472_ _5215_/A _4399_/B _5472_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_129_196 VGND VPWR sky130_fd_sc_hd__decap_12
X_7211_ _7615_/Q la_data_in[109] _7147_/X _7211_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_4423_ _4291_/A _4903_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_144_166 VGND VPWR sky130_fd_sc_hd__decap_12
X_7142_ _7616_/Q _7142_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_193_1160 VGND VPWR sky130_fd_sc_hd__decap_12
X_4354_ _4301_/A _4301_/B _4301_/X _4368_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_141_840 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_754 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_787 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_1038 VGND VPWR sky130_fd_sc_hd__decap_12
X_7073_ _7619_/Q _7073_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_154_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_798 VGND VPWR sky130_fd_sc_hd__decap_12
X_4285_ _4283_/X _4284_/X _4283_/X _4284_/X _4285_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_150_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_895 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_426 VGND VPWR sky130_fd_sc_hd__decap_12
X_6024_ _5051_/Y _6148_/A _6023_/X _6024_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_86_459 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_971 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_323 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_654 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_518 VGND VPWR sky130_fd_sc_hd__fill_1
X_6926_ _7648_/Q _6926_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_3229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_800 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6857_ _6857_/A _6857_/B _6857_/X VGND VPWR sky130_fd_sc_hd__and2_4
XPHY_2539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5808_ _5805_/X _5806_/X _5805_/X _5806_/X _5808_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_10_404 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_940 VGND VPWR sky130_fd_sc_hd__decap_12
X_6788_ _7676_/Q la_data_in[42] _6723_/X _6788_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XPHY_1849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_1101 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_578 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_448 VGND VPWR sky130_fd_sc_hd__decap_8
X_5739_ _5736_/X _5737_/X _5749_/A _5739_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_164_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_601 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_954 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_740 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_807 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1093 VGND VPWR sky130_fd_sc_hd__decap_12
X_7409_ io_oeb[4] _7409_/LO VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_136_678 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_497 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1203 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_1211 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_575 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_908 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_993 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_857 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_98 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_367 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1048 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_851 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_63 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_4475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_581 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_220 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_361 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_562 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_534 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1005 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_475 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_935 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_328 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_394 VGND VPWR sky130_fd_sc_hd__decap_3
X_4070_ _4070_/A _4070_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_95_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1060 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_407 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_443 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_301 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_1123 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_632 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1047 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_654 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_345 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_498 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1126 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_1069 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_816 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_304 VGND VPWR sky130_fd_sc_hd__fill_1
X_7760_ _6259_/X _5507_/A _7797_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4972_ _4932_/X _4933_/X _4922_/X _4934_/X _4972_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_6711_ _6709_/Y _6710_/Y _6709_/Y _6710_/Y _6770_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_3923_ _4218_/B _3949_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_211_118 VGND VPWR sky130_fd_sc_hd__decap_6
X_7691_ _6683_/X _6615_/A _7696_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_177_501 VGND VPWR sky130_fd_sc_hd__decap_4
X_6642_ _6639_/Y _6640_/Y _6639_/Y _6640_/Y _6642_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_3854_ _4716_/A _5137_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_20_735 VGND VPWR sky130_fd_sc_hd__decap_8
X_6573_ _6548_/X _6571_/X _6572_/X _6573_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_146_910 VGND VPWR sky130_fd_sc_hd__decap_12
X_3785_ _7808_/Q _3786_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_164_239 VGND VPWR sky130_fd_sc_hd__decap_12
X_5524_ _5319_/X _5320_/X _5318_/X _5321_/X _5524_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_195_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_678 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_464 VGND VPWR sky130_fd_sc_hd__decap_12
X_5455_ _5399_/X _5452_/X _5453_/X _5454_/X _5455_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_105_306 VGND VPWR sky130_fd_sc_hd__decap_8
X_4406_ _4919_/A _4460_/B _4408_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_114_840 VGND VPWR sky130_fd_sc_hd__decap_12
X_5386_ _5375_/X _5376_/X _5374_/X _5377_/X _5386_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_7125_ _7084_/X _7124_/X _7114_/X _7125_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_4337_ _4336_/A _4335_/X _4336_/X _4337_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_141_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_501 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_724 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1016 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_448 VGND VPWR sky130_fd_sc_hd__decap_12
X_7056_ la_data_in[87] _7057_/B VGND VPWR sky130_fd_sc_hd__inv_8
X_4268_ _4847_/A _4399_/B _4268_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_41_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_971 VGND VPWR sky130_fd_sc_hd__fill_1
X_6007_ _5459_/X _5518_/Y _6006_/X _6008_/B VGND VPWR sky130_fd_sc_hd__o21ai_4
X_4199_ _4155_/X _4196_/X _4197_/Y _4198_/X _4200_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_83_930 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_367 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_687 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_827 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_495 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_197 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6909_ _6869_/X _6908_/X _6905_/X _6909_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XPHY_2325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_129 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_512 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_44 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_652 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_342 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_88 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_757 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_717 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_526 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_656 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_570 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_486 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_626 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_41 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1003 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_990 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_372 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_735 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1063 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_854 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_908 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_705 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_356 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_602 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1160 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_1171 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_849 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1121 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_523 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_692 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_167 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1192 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1187 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_921 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_954 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_750 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_946 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_497 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_142_434 VGND VPWR sky130_fd_sc_hd__decap_12
X_5240_ _3846_/X _4459_/B _5240_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_46_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1130 VGND VPWR sky130_fd_sc_hd__fill_1
X_5171_ _5171_/A _4455_/B _5172_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_69_746 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1008 VGND VPWR sky130_fd_sc_hd__fill_1
X_4122_ _4494_/A _4122_/B _4122_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_151_1125 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_919 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_727 VGND VPWR sky130_fd_sc_hd__decap_12
X_4053_ _7740_/Q _4054_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_65_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_922 VGND VPWR sky130_fd_sc_hd__decap_3
X_7812_ _3761_/Y _7812_/Q _7810_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_24_315 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_1054 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_186 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_27 VGND VPWR sky130_fd_sc_hd__decap_12
X_7743_ _6336_/Y _7743_/Q _7806_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4955_ _4914_/X _4920_/X _4913_/X _4921_/X _4955_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_75_1251 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_117 VGND VPWR sky130_fd_sc_hd__decap_12
X_3906_ wbs_dat_i[0] _3882_/X _3907_/C VGND VPWR sky130_fd_sc_hd__nor2_4
X_7674_ _6795_/X _6727_/A _7756_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_20_510 VGND VPWR sky130_fd_sc_hd__decap_8
X_4886_ _4886_/A _4888_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_20_532 VGND VPWR sky130_fd_sc_hd__decap_12
X_6625_ la_data_in[22] _6625_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_178_898 VGND VPWR sky130_fd_sc_hd__decap_12
X_3837_ _3757_/A _3838_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_192_312 VGND VPWR sky130_fd_sc_hd__decap_12
X_6556_ la_data_in[15] _6556_/B _6556_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_3768_ wbs_dat_i[17] _3790_/B _3768_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_193_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_913 VGND VPWR sky130_fd_sc_hd__decap_12
X_5507_ _5507_/A _5445_/Y _5507_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_3_208 VGND VPWR sky130_fd_sc_hd__decap_12
X_6487_ _6487_/A _6487_/B _6487_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_3699_ wbs_adr_i[9] wbs_adr_i[8] wbs_adr_i[11] wbs_adr_i[10] _3699_/X VGND VPWR sky130_fd_sc_hd__or4_4
X_5438_ _5434_/X _5437_/X _5434_/X _5437_/X _5438_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_105_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1069 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_489 VGND VPWR sky130_fd_sc_hd__decap_12
X_5369_ _5366_/X _5367_/X _5368_/X _5371_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_126_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_681 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1266 VGND VPWR sky130_fd_sc_hd__decap_8
X_7108_ _7092_/X _7107_/X _7024_/X _7108_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_59_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_727 VGND VPWR sky130_fd_sc_hd__decap_4
X_7039_ _7037_/Y _7038_/Y _7039_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_102_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_941 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_963 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_440 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_906 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_782 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_473 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_175 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_849 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_326 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_629 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_145 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_98 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_487 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_381 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_673 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1048 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_554 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_239 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_97 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_902 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_453 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1212 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_581 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1245 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_253 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_467 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_264 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_938 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1240 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_952 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_733 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_202_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1126 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_1069 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_112 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1268 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_679 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_318 VGND VPWR sky130_fd_sc_hd__decap_12
X_4740_ _4716_/X _4720_/X _4716_/X _4720_/X _4740_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_3390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_684 VGND VPWR sky130_fd_sc_hd__decap_12
X_4671_ _4624_/X _4629_/X _4624_/X _4629_/X _4671_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_159_386 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_312 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_1003 VGND VPWR sky130_fd_sc_hd__decap_12
X_6410_ la_data_in[117] _6410_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_174_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_548 VGND VPWR sky130_fd_sc_hd__fill_1
X_7390_ io_in[32] _7390_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_175_879 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_902 VGND VPWR sky130_fd_sc_hd__fill_1
X_6341_ _4122_/B _6348_/B _6343_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_192_1203 VGND VPWR sky130_fd_sc_hd__decap_12
X_6272_ _6269_/Y _6270_/X _6273_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_143_787 VGND VPWR sky130_fd_sc_hd__decap_6
X_5223_ _5213_/X _5220_/X _5221_/X _5222_/X _5223_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_115_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1020 VGND VPWR sky130_fd_sc_hd__decap_12
X_5154_ _5143_/X _5147_/X _5146_/X _5154_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_9_1155 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_885 VGND VPWR sky130_fd_sc_hd__decap_8
X_4105_ _4104_/A _4104_/B _4104_/Y _6095_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_111_684 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_5085_ _5171_/A _4597_/B _5087_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_116_1097 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_80 VGND VPWR sky130_fd_sc_hd__fill_1
X_4036_ _4036_/A _4036_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_112_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_410 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_741 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_107 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_977 VGND VPWR sky130_fd_sc_hd__decap_12
X_5987_ _5884_/X _5908_/X _5909_/X _5986_/X _6280_/A VGND VPWR sky130_fd_sc_hd__o22a_4
XPHY_118 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_605 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_129 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_178 VGND VPWR sky130_fd_sc_hd__decap_12
X_4938_ _4912_/X _4937_/X _4912_/X _4937_/X _4938_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7726_ _6457_/X _7726_/Q _7785_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_75_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1043 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_830 VGND VPWR sky130_fd_sc_hd__decap_12
X_4869_ _4652_/X _4660_/X _4644_/X _4661_/X _4869_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_7657_ _6907_/X _6840_/A _7707_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_166_846 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_373 VGND VPWR sky130_fd_sc_hd__decap_3
X_6608_ _6606_/Y _6608_/B _6608_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_7588_ _7588_/HI la_data_out[115] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_123_1079 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_838 VGND VPWR sky130_fd_sc_hd__decap_12
X_6539_ _6524_/X _6539_/B _6539_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_21_56 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_957 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_434 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_745 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_1183 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1025 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_727 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1039 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_53 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_123 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_9 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_752 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_426 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_476 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1121 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_148 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_684 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_846 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1138 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1206 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_384 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_849 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_765 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_916 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_550 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_787 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_746 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1212 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_800 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_1158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_1010 VGND VPWR sky130_fd_sc_hd__decap_12
X_5910_ _5906_/X _5907_/X _5906_/X _5907_/X _5910_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_410 VGND VPWR sky130_fd_sc_hd__decap_4
X_6890_ _6878_/X _6888_/X _6889_/Y _6890_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_207_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1062 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_752 VGND VPWR sky130_fd_sc_hd__decap_8
X_5841_ _5824_/X _5840_/X _5841_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_35_977 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_605 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_925 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_706 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_947 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_638 VGND VPWR sky130_fd_sc_hd__decap_3
X_5772_ _5768_/X _5769_/X _5770_/X _5771_/X _5772_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_4723_ _4715_/X _4721_/X _4715_/X _4721_/X _4723_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7511_ _7511_/HI la_data_out[38] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_72_1265 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_159 VGND VPWR sky130_fd_sc_hd__decap_3
X_7442_ io_oeb[37] _7442_/LO VGND VPWR sky130_fd_sc_hd__conb_1
X_4654_ _4654_/A _4666_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_30_693 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_710 VGND VPWR sky130_fd_sc_hd__decap_12
X_7373_ _5534_/Y _7355_/X _7372_/X wbs_dat_o[20] VGND VPWR sky130_fd_sc_hd__o21ai_4
X_4585_ _4580_/Y _4584_/X _4580_/Y _4584_/X _4585_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_128_581 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_337 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_1276 VGND VPWR sky130_fd_sc_hd__fill_1
X_6324_ _6340_/A _6334_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_162_359 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_754 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_679 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_798 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_415 VGND VPWR sky130_fd_sc_hd__decap_12
X_6255_ _6255_/A _6255_/B _7761_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_192_1066 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_59 VGND VPWR sky130_fd_sc_hd__fill_2
X_5206_ _5197_/X _5203_/X _5204_/X _5205_/X _5206_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_6186_ _4806_/A _4806_/B _6150_/B _6186_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_112_971 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_351 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_513 VGND VPWR sky130_fd_sc_hd__decap_12
X_5137_ _5137_/A _4852_/B _5137_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_85_855 VGND VPWR sky130_fd_sc_hd__fill_1
X_5068_ _5066_/X _5067_/X _5065_/X _5068_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XPHY_4805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_771 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_922 VGND VPWR sky130_fd_sc_hd__decap_4
X_4019_ _4399_/B _4122_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_84_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1121 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_281 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_251 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_129_1255 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1029 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_89 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1119 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_200_227 VGND VPWR sky130_fd_sc_hd__decap_12
X_7709_ _7709_/D _6501_/A _7658_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_32_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_849 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_551 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1242 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_175_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1109 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_531 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_839 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1013 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_313 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_741 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_936 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1219 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_446 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_468 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_693 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_642 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1025 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_624 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_1047 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_196 VGND VPWR sky130_fd_sc_hd__decap_12
X_4370_ _3689_/A _4295_/A _4189_/A _4293_/X _4370_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_125_562 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_947 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_881 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_180_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_757 VGND VPWR sky130_fd_sc_hd__decap_12
X_6040_ _6070_/A _6139_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_3_391 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_576 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1192 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_708 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_803 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_376 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_398 VGND VPWR sky130_fd_sc_hd__decap_12
X_6942_ la_data_in[73] _6942_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_47_590 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_379 VGND VPWR sky130_fd_sc_hd__decap_12
X_6873_ _6837_/Y _6838_/Y _6872_/X _6873_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_179_245 VGND VPWR sky130_fd_sc_hd__decap_12
X_5824_ _3904_/X _4346_/B _5824_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_194_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_5755_ _5754_/A _5710_/Y _5754_/X _5755_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_210_547 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_654 VGND VPWR sky130_fd_sc_hd__decap_12
X_4706_ _4693_/X _4703_/X _4704_/X _4705_/X _4706_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_175_440 VGND VPWR sky130_fd_sc_hd__decap_12
X_5686_ _5681_/X _5685_/X _5684_/X _5686_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_176_996 VGND VPWR sky130_fd_sc_hd__decap_8
X_4637_ _4630_/X _4636_/X _4630_/X _4636_/X _4637_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7425_ io_oeb[20] _7425_/LO VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_163_635 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_410 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1049 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_977 VGND VPWR sky130_fd_sc_hd__decap_4
X_4568_ _4568_/A _4512_/B _4568_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7356_ io_in[22] _7356_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_162_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_318 VGND VPWR sky130_fd_sc_hd__decap_12
X_6307_ _3733_/A _6306_/Y _7749_/D VGND VPWR sky130_fd_sc_hd__nor2_4
X_7287_ io_in[10] _7288_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_4499_ _4499_/A _4570_/B _4500_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_6238_ _6198_/A _6238_/B _6240_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_103_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_6169_ _5003_/Y _6158_/X _6144_/X _6169_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_134_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_844 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_663 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_354 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_56 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_88 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_379 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_796 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_21 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_947 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_284 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_727 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_587 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_1096 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_428 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_1017 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_952 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_963 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_805 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_451 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_760 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_816 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_827 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_315 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_944 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1209 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_623 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_562 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_166 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_1001 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_177 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_59 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1094 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1097 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_874 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_1067 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_350 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_110_738 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_647 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_658 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_825 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1062 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1099 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_1043 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1046 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_593 VGND VPWR sky130_fd_sc_hd__decap_8
X_3870_ _4718_/A _5348_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_56_1057 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_407 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1038 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_749 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_290 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_940 VGND VPWR sky130_fd_sc_hd__decap_12
X_5540_ _5536_/X _5539_/X _5536_/X _5539_/X _5540_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_157_440 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_974 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_450 VGND VPWR sky130_fd_sc_hd__decap_8
X_5471_ _5466_/X _5470_/X _5469_/X _5471_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_8_494 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_443 VGND VPWR sky130_fd_sc_hd__decap_12
X_4422_ _3720_/A _4569_/B _4422_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7210_ _7210_/A _7203_/X _7209_/Y _7210_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_173_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_178 VGND VPWR sky130_fd_sc_hd__decap_12
X_7141_ _7210_/A _7077_/A _7140_/X _7141_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_119_1210 VGND VPWR sky130_fd_sc_hd__decap_8
X_4353_ _4326_/X _4341_/X _4351_/X _4352_/X _4353_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_99_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1126 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_852 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_906 VGND VPWR sky130_fd_sc_hd__decap_8
X_7072_ _7070_/Y _7071_/Y _7072_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_87_928 VGND VPWR sky130_fd_sc_hd__decap_8
X_4284_ _4237_/X _4238_/X _4237_/X _4238_/X _4284_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_373 VGND VPWR sky130_fd_sc_hd__decap_12
X_6023_ _5051_/Y _6011_/X _6017_/Y _6022_/X _6023_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_100_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_438 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_641 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_663 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_696 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_318 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_666 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6925_ _6923_/A _6922_/A _6924_/X _7650_/D VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_70_828 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_711 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_733 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1263 VGND VPWR sky130_fd_sc_hd__decap_12
X_6856_ la_data_in[50] _6857_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_168_716 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_300 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_541 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_906 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5807_ _5807_/A _5807_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_1828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_928 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3999_ _3999_/A _4000_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_6787_ _6766_/X _6784_/X _6786_/Y _7677_/D VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_149_952 VGND VPWR sky130_fd_sc_hd__decap_3
X_5738_ _5736_/X _5737_/X _5749_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_164_922 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_613 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_827 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1061 VGND VPWR sky130_fd_sc_hd__decap_6
X_5669_ _5656_/X _5657_/X _5658_/X _5669_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_135_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_337 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_966 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_752 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_7408_ io_oeb[3] _7408_/LO VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_124_819 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_103 VGND VPWR sky130_fd_sc_hd__decap_8
X_7339_ io_in[19] _7340_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_1_114 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_532 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1237 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_395 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_760 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_611 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_313 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_869 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_20 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1027 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_379 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1013 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_812 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_593 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_232 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_373 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_215 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_546 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_900 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_782 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_410 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1112 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_752 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1156 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_487 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_947 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_1_0_wb_clk_i clkbuf_1_0_1_wb_clk_i/X clkbuf_2_1_1_wb_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_141_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_928 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_362 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_180 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_419 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1139 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1059 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_975 VGND VPWR sky130_fd_sc_hd__decap_12
X_4971_ _4967_/X _4970_/X _4967_/X _4970_/X _4971_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_149_1269 VGND VPWR sky130_fd_sc_hd__decap_8
X_6710_ la_data_in[46] _6710_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_3922_ _4394_/B _4218_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_205_672 VGND VPWR sky130_fd_sc_hd__decap_12
X_7690_ _7690_/D _7690_/Q _7696_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_60_861 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_703 VGND VPWR sky130_fd_sc_hd__decap_12
X_3853_ _5171_/A _4716_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_6641_ _6641_/A la_data_in[16] _6705_/A VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_165_708 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_259 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1130 VGND VPWR sky130_fd_sc_hd__decap_3
X_3784_ _3743_/A _3791_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_6572_ _6670_/A _6572_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_121_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_922 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_624 VGND VPWR sky130_fd_sc_hd__decap_12
X_5523_ _4765_/X _4766_/X _4765_/X _4766_/X _5523_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_69_1204 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_123 VGND VPWR sky130_fd_sc_hd__decap_12
X_5454_ _5399_/X _5452_/X _5399_/X _5452_/X _5454_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_195_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_785 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_476 VGND VPWR sky130_fd_sc_hd__decap_12
X_4405_ _4391_/X _4397_/X _4403_/X _4404_/X _4405_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_5385_ _5381_/X _5382_/X _5383_/Y _5384_/X _5385_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_126_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_852 VGND VPWR sky130_fd_sc_hd__decap_6
X_4336_ _4336_/A _4335_/X _4336_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7124_ _7058_/A la_data_in[86] _7060_/X _7124_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_115_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1028 VGND VPWR sky130_fd_sc_hd__decap_12
X_7055_ _7055_/A _7057_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_4267_ _4498_/A _4925_/B _4269_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_115_59 VGND VPWR sky130_fd_sc_hd__fill_2
X_6006_ _6006_/A _6006_/B _6006_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_132_1240 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1183 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_151 VGND VPWR sky130_fd_sc_hd__decap_12
X_4198_ _4155_/X _4196_/X _4155_/X _4196_/X _4198_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_55_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_847 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_942 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_666 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_3005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_305 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_379 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_699 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_839 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_159 VGND VPWR sky130_fd_sc_hd__decap_12
X_6908_ _6843_/A la_data_in[54] _6845_/X _6908_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XPHY_3049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_563 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6839_ _6837_/Y _6838_/Y _6837_/Y _6838_/Y _6872_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_1625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_664 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_585 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_141 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_354 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1088 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1252 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_246 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_729 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_538 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_1274 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_944 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_668 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_424 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_498 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_638 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_423 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1061 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_863 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1151 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_467 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_811 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_53 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1015 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_384 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_747 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_866 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_877 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_961 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_27 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_791 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_313 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_666 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_463 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_368 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1183 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_4262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1021 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_179 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_894 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_1098 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_888 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_966 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_733 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_958 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_294 VGND VPWR sky130_fd_sc_hd__decap_8
X_5170_ _4749_/A _4748_/B _5172_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_68_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_4121_ _4113_/X _4120_/X _4113_/X _4120_/X _4121_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_321 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_758 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1137 VGND VPWR sky130_fd_sc_hd__decap_12
X_4052_ _4049_/X _4050_/X _4051_/X _4059_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_84_739 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_964 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1022 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_761 VGND VPWR sky130_fd_sc_hd__fill_2
X_7811_ _3769_/Y _7811_/Q _7774_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_188_1082 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_783 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_1066 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_956 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_293 VGND VPWR sky130_fd_sc_hd__decap_12
X_7742_ _6339_/Y _3999_/A _7810_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_178_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_349 VGND VPWR sky130_fd_sc_hd__fill_2
X_4954_ _4907_/X _4908_/X _4900_/X _4909_/X _4954_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_149_1099 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_809 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1211 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_196_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_3905_ _3904_/X _3897_/B _3907_/B VGND VPWR sky130_fd_sc_hd__and2_4
X_7673_ _6798_/X _7673_/Q _7758_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4885_ _4819_/X _4836_/X _4818_/X _4837_/X _4885_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_6624_ _6624_/A _6624_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_119_900 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_544 VGND VPWR sky130_fd_sc_hd__decap_12
X_3836_ _4678_/A _5420_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_192_324 VGND VPWR sky130_fd_sc_hd__decap_12
X_3767_ _5058_/A _3767_/B _3767_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_6555_ io_out[0] _6554_/X _6556_/B VGND VPWR sky130_fd_sc_hd__xnor2_4
XFILLER_69_1001 VGND VPWR sky130_fd_sc_hd__decap_4
X_5506_ _5495_/X _5496_/X _5494_/X _5497_/X _5506_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_134_925 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_999 VGND VPWR sky130_fd_sc_hd__decap_12
X_3698_ wbs_adr_i[13] wbs_adr_i[12] wbs_adr_i[15] wbs_adr_i[14] _3700_/A VGND VPWR
+ sky130_fd_sc_hd__or4_4
X_6486_ _6426_/X _6484_/X _6485_/Y _6486_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_161_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1064 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_947 VGND VPWR sky130_fd_sc_hd__decap_12
X_5437_ _5435_/X _5436_/X _5435_/X _5436_/X _5437_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_105_159 VGND VPWR sky130_fd_sc_hd__decap_12
X_5368_ _5366_/X _5367_/X _5368_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_160_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_693 VGND VPWR sky130_fd_sc_hd__decap_8
X_7107_ _7040_/A la_data_in[92] _7042_/X _7107_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_43_1218 VGND VPWR sky130_fd_sc_hd__fill_2
X_4319_ _4253_/A _4318_/X _4253_/A _4318_/X _4320_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_5299_ _5133_/X _5134_/X _5127_/X _5135_/X _5299_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_206_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_257 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_354 VGND VPWR sky130_fd_sc_hd__decap_12
X_7038_ la_data_in[93] _7038_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_59_279 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_633 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_986 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_485 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_918 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_33 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1188 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_428 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1130 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_989 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_861 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_499 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_371 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_190 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_685 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_184 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_869 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1112 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_379 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_465 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1137 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_231 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_242 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_660 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_253 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_264 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_511 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_544 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_216 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_1212 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1121 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1252 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_603 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_756 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1108 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_293 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_135 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_157 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_940 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1072 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_814 VGND VPWR sky130_fd_sc_hd__fill_1
X_4670_ _4665_/X _4669_/X _4668_/X _4670_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_202_483 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_696 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_159_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_886 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_1015 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1111 VGND VPWR sky130_fd_sc_hd__decap_12
X_6340_ _6340_/A _6348_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_143_733 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_581 VGND VPWR sky130_fd_sc_hd__decap_8
X_6271_ _6269_/Y _6270_/X _6273_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_192_1215 VGND VPWR sky130_fd_sc_hd__decap_12
X_5222_ _5213_/X _5220_/X _5213_/X _5220_/X _5222_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_142_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1062 VGND VPWR sky130_fd_sc_hd__decap_12
X_5153_ _5121_/X _5152_/X _5121_/X _5152_/X _5153_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_116_1032 VGND VPWR sky130_fd_sc_hd__fill_2
X_4104_ _4104_/A _4104_/B _4104_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_5084_ _5420_/A _4595_/B _5084_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_56_205 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_536 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_227 VGND VPWR sky130_fd_sc_hd__decap_6
X_4035_ _4035_/A _4036_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_186_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_750 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_794 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_647 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_753 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_108 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_764 VGND VPWR sky130_fd_sc_hd__decap_8
X_5986_ _5910_/X _5926_/X _5985_/X _5986_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XPHY_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_617 VGND VPWR sky130_fd_sc_hd__decap_12
X_7725_ _7725_/D _7725_/Q _7785_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4937_ _4935_/X _4936_/X _4935_/X _4936_/X _4937_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_75_1093 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_127_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_842 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_20 _5383_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_7656_ _6910_/X _6843_/A _7707_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_193_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_864 VGND VPWR sky130_fd_sc_hd__decap_12
X_4868_ _4859_/X _4867_/X _4859_/X _4867_/X _4868_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_138_527 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1036 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_165_313 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_184 VGND VPWR sky130_fd_sc_hd__decap_12
X_6607_ la_data_in[28] _6608_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_166_858 VGND VPWR sky130_fd_sc_hd__decap_12
X_3819_ _4547_/A _4653_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_7587_ _7587_/HI la_data_out[114] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_181_806 VGND VPWR sky130_fd_sc_hd__decap_6
X_4799_ _4797_/X _4798_/X _4797_/X _4798_/X _4799_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_20_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_251 VGND VPWR sky130_fd_sc_hd__decap_12
X_6538_ _6527_/A _6526_/Y _6527_/X _6537_/X _6539_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_134_711 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_880 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_936 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_969 VGND VPWR sky130_fd_sc_hd__decap_6
X_6469_ _7721_/Q la_data_in[119] _6405_/X _6469_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_133_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_906 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_574 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_788 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1195 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_739 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1217 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_709 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_964 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_65 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_400 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_135 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_438 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1242 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_641 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_269 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_910 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_516 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_330 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_302 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_1008 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_280 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_886 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_363 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_15 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_335 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1218 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_666 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_396 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_733 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_390 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_758 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_1232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_471 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_227 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_249 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_901 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1022 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_783 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_794 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_179_405 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_586 VGND VPWR sky130_fd_sc_hd__decap_12
X_5840_ _5825_/X _5839_/B _5839_/X _5840_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_185_1074 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1099 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_937 VGND VPWR sky130_fd_sc_hd__decap_8
X_5771_ _5768_/X _5769_/X _5768_/X _5769_/X _5771_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_803 VGND VPWR sky130_fd_sc_hd__fill_1
X_7510_ _7510_/HI la_data_out[37] VGND VPWR sky130_fd_sc_hd__conb_1
X_4722_ _4452_/X _4457_/X _4452_/X _4457_/X _4722_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_175_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_847 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_184 VGND VPWR sky130_fd_sc_hd__decap_12
X_7441_ io_oeb[36] _7441_/LO VGND VPWR sky130_fd_sc_hd__conb_1
X_4653_ _4653_/A _4653_/B _4653_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_163_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_508 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_305 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_560 VGND VPWR sky130_fd_sc_hd__decap_12
X_7372_ _3738_/X _7370_/X _7371_/Y _7364_/X _7372_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_4584_ _4581_/X _4583_/X _4581_/X _4583_/X _4584_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_116_722 VGND VPWR sky130_fd_sc_hd__fill_2
X_6323_ _6323_/A _7264_/B _6340_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_196_1170 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1004 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_541 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1154 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_192_1034 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_574 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_788 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_6254_ _5383_/Y _6091_/X _6190_/X _6255_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_130_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1176 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1149 VGND VPWR sky130_fd_sc_hd__decap_8
X_5205_ _5197_/X _5203_/X _5197_/X _5203_/X _5205_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6185_ _6185_/A _6185_/B _7772_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_69_363 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_983 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_672 VGND VPWR sky130_fd_sc_hd__decap_6
X_5136_ _5127_/X _5135_/X _5127_/X _5135_/X _5136_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_84_300 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_205 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_385 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_525 VGND VPWR sky130_fd_sc_hd__decap_12
X_5067_ _4512_/A _4493_/X _5067_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_123_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4018_ _4748_/B _4399_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_783 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1133 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1136 VGND VPWR sky130_fd_sc_hd__fill_1
X_5969_ _5967_/X _5968_/X _5969_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_179_961 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_408 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1111 VGND VPWR sky130_fd_sc_hd__decap_12
X_7708_ _6574_/X _7708_/Q _7707_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_200_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_56 VGND VPWR sky130_fd_sc_hd__decap_12
X_7639_ _7020_/X _7639_/Q _7624_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_194_975 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_182 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_563 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1257 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_736 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_543 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_257 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_565 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1025 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1154 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_325 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_794 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_714 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_753 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_550 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_556 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_477 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_959 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_611 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_964 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_441 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_131 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_154 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_997 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1059 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_714 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_893 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1032 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1098 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_815 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_388 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_528 VGND VPWR sky130_fd_sc_hd__decap_12
X_6941_ _7643_/Q _6941_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_93_196 VGND VPWR sky130_fd_sc_hd__decap_12
X_6872_ _6872_/A _6871_/X _6872_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_23_904 VGND VPWR sky130_fd_sc_hd__decap_8
X_5823_ _5812_/X _5813_/X _5812_/X _5813_/X _5823_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_179_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_706 VGND VPWR sky130_fd_sc_hd__fill_1
X_5754_ _5754_/A _5710_/Y _5754_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_194_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_559 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1142 VGND VPWR sky130_fd_sc_hd__decap_3
X_4705_ _4693_/X _4703_/X _4693_/X _4703_/X _4705_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_33_1036 VGND VPWR sky130_fd_sc_hd__fill_1
X_5685_ _5684_/A _5684_/B _5684_/X _5685_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_175_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_666 VGND VPWR sky130_fd_sc_hd__decap_12
X_7424_ io_oeb[19] _7424_/LO VGND VPWR sky130_fd_sc_hd__conb_1
X_4636_ _4631_/X _4635_/X _4631_/X _4635_/X _4636_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_194_1107 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_7355_ _7354_/X _7355_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_163_669 VGND VPWR sky130_fd_sc_hd__fill_2
X_4567_ _4566_/A _4565_/X _4581_/B _4567_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_144_861 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_703 VGND VPWR sky130_fd_sc_hd__decap_8
X_6306_ _5978_/B _6073_/X _6305_/X _7749_/Q _6084_/X _6306_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_144_894 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_511 VGND VPWR sky130_fd_sc_hd__decap_12
X_7286_ _4070_/A _7260_/B _7286_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_4498_ _4498_/A _4498_/B _4500_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_171_691 VGND VPWR sky130_fd_sc_hd__decap_4
X_6237_ _6197_/X _6198_/B _5518_/A _6238_/B VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_170_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_257 VGND VPWR sky130_fd_sc_hd__decap_12
X_6168_ _6165_/Y _6166_/X _6319_/C _6168_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_97_480 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_856 VGND VPWR sky130_fd_sc_hd__decap_12
X_5119_ _5071_/X _5118_/X _5071_/X _5118_/X _5119_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_85_653 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_141 VGND VPWR sky130_fd_sc_hd__decap_12
X_6099_ _6095_/Y _6098_/Y _4104_/Y _6099_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_27_23 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1228 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_826 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_208 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_68 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_3_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A clkbuf_4_7_0_wb_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_4669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_403 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_33 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_959 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_739 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_611 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_1212 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1242 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_1029 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_986 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_839 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_327 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_349 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_390 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_189 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_841 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_300 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_631 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_322 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_867 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_810 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_712 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_189_566 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1055 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_419 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_931 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_110 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_280 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_291 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_463 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_581 VGND VPWR sky130_fd_sc_hd__decap_12
X_5470_ _5467_/X _5468_/X _5469_/X _5470_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_172_411 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_484 VGND VPWR sky130_fd_sc_hd__fill_1
X_4421_ _4360_/X _4366_/X _4360_/X _4366_/X _4430_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_172_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_989 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_712 VGND VPWR sky130_fd_sc_hd__decap_3
X_7140_ _7618_/Q la_data_in[80] _7140_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_160_639 VGND VPWR sky130_fd_sc_hd__fill_2
X_4352_ _4326_/X _4341_/X _4326_/X _4341_/X _4352_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_113_511 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1105 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_745 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_190 VGND VPWR sky130_fd_sc_hd__decap_12
X_4283_ _4270_/X _4271_/X _4269_/X _4283_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_7071_ la_data_in[82] _7071_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_6022_ _6018_/X _5030_/Y _5014_/X _6021_/Y _6022_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_98_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_995 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_196 VGND VPWR sky130_fd_sc_hd__fill_1
X_6924_ _6860_/A la_data_in[48] _6924_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_3209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_678 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_550 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_120_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_723 VGND VPWR sky130_fd_sc_hd__decap_8
X_6855_ _7652_/Q _6857_/A VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_2519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1253 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1275 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_728 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_312 VGND VPWR sky130_fd_sc_hd__fill_2
X_5806_ _5420_/A _5294_/B _5806_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_1818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_553 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_525 VGND VPWR sky130_fd_sc_hd__decap_12
X_6786_ _6766_/X _6784_/X _6785_/X _6786_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XPHY_1829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3998_ _3971_/X _3982_/Y _4027_/B _3998_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_210_345 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_597 VGND VPWR sky130_fd_sc_hd__fill_1
X_5737_ _3850_/Y _4820_/B _5737_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_200_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_806 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_839 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1002 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_934 VGND VPWR sky130_fd_sc_hd__decap_12
X_5668_ _5668_/A _5667_/X _5668_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_191_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_293 VGND VPWR sky130_fd_sc_hd__decap_12
X_7407_ io_oeb[2] _7407_/LO VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_135_135 VGND VPWR sky130_fd_sc_hd__decap_12
X_4619_ _4617_/X _4618_/X _4617_/X _4618_/X _4619_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_164_978 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_764 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_1210 VGND VPWR sky130_fd_sc_hd__decap_8
X_5599_ _4548_/A _5123_/B _5599_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_85_1221 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_7338_ _7338_/A _7321_/B _7338_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_116_371 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_649 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_126 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_907 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_137 VGND VPWR sky130_fd_sc_hd__decap_8
X_7269_ _7779_/Q _7260_/B _7269_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_132_875 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_341 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1249 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_588 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_951 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1090 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_130 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_472 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_837 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_1036 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_634 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_325 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_173_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_196 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_818 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_166 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_734 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1025 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_391 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1258 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_385 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_879 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_186_558 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_912 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_923 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1124 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_499 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_831 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_374 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1221 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1013 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_686 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_111 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1106 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_987 VGND VPWR sky130_fd_sc_hd__decap_12
X_4970_ _4968_/X _4969_/X _4968_/X _4969_/X _4970_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_52_829 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_306 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_550 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_317 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_330 VGND VPWR sky130_fd_sc_hd__decap_12
X_3921_ _4743_/B _4394_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_32_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_684 VGND VPWR sky130_fd_sc_hd__decap_12
X_6640_ la_data_in[17] _6640_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_3852_ _4680_/A _5171_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_60_873 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_715 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_249 VGND VPWR sky130_fd_sc_hd__fill_1
X_6571_ _7708_/Q la_data_in[10] _6506_/X _6571_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_34_1142 VGND VPWR sky130_fd_sc_hd__decap_12
X_3783_ _3769_/A _3781_/X _3782_/Y _3783_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_192_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1123 VGND VPWR sky130_fd_sc_hd__decap_12
X_5522_ _4789_/X _4790_/X _4789_/X _4790_/X _5522_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_934 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_636 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_1216 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_135 VGND VPWR sky130_fd_sc_hd__decap_12
X_5453_ _5447_/X _5448_/X _5446_/Y _5449_/X _5453_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_172_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_4404_ _4391_/X _4397_/X _4391_/X _4397_/X _4404_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_520 VGND VPWR sky130_fd_sc_hd__decap_12
X_5384_ _5381_/X _5382_/X _5381_/X _5382_/X _5384_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7123_ _7085_/X _7121_/X _7122_/Y _7123_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_113_330 VGND VPWR sky130_fd_sc_hd__decap_4
X_4335_ _4570_/A _4590_/B _4335_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_114_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_428 VGND VPWR sky130_fd_sc_hd__fill_1
X_7054_ _7052_/Y _7053_/Y _7052_/Y _7053_/Y _7119_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_119_1096 VGND VPWR sky130_fd_sc_hd__fill_2
X_4266_ _4260_/X _4265_/X _4264_/X _4266_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_6005_ _6005_/A _6005_/B _5332_/X _6005_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_132_1252 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_815 VGND VPWR sky130_fd_sc_hd__decap_8
X_4197_ _7780_/Q _4197_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_95_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_163 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_837 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_859 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_954 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_196 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_166 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_317 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6907_ _6870_/X _6904_/X _6906_/Y _6907_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XPHY_3039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_621 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6838_ la_data_in[56] _6838_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_1604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_361 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1067 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_597 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_676 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6769_ _6712_/Y _6714_/B _6714_/X _6768_/X _6769_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XPHY_1659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_956 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_753 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_56 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_764 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_477 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1073 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_759 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_973 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_932 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_325 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_86 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_306 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_520 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_4274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_503 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_812 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1033 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_531 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_672 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_300 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_654 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_74 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_558 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_867 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_74 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_934 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_7 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_978 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_778 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1108 VGND VPWR sky130_fd_sc_hd__decap_12
X_4120_ _4118_/X _4119_/X _4117_/X _4120_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_96_534 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1179 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_1149 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_1269 VGND VPWR sky130_fd_sc_hd__decap_8
X_4051_ _4049_/X _4050_/X _4051_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_96_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_366 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_623 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_740 VGND VPWR sky130_fd_sc_hd__fill_2
X_7810_ _3776_/Y _7810_/Q _7810_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_25_818 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1034 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_1094 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_795 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_328 VGND VPWR sky130_fd_sc_hd__decap_8
X_7741_ _6343_/Y _7741_/Q _7806_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_206_971 VGND VPWR sky130_fd_sc_hd__decap_12
X_4953_ _4951_/X _4952_/B _4952_/X _4953_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_80_968 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_380 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_812 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1215 VGND VPWR sky130_fd_sc_hd__decap_12
X_3904_ _5215_/A _3904_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_7672_ _6801_/X _7672_/Q _7756_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_189_171 VGND VPWR sky130_fd_sc_hd__decap_12
X_4884_ _4881_/A _4880_/X _4883_/X _4884_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_60_670 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_361 VGND VPWR sky130_fd_sc_hd__decap_12
X_6623_ _6621_/Y _6623_/B _6623_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_3835_ _4455_/A _4678_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_137_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_912 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_556 VGND VPWR sky130_fd_sc_hd__decap_12
X_6554_ _6492_/Y _6493_/Y _6553_/X _6554_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_3766_ _4503_/A _5058_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_146_742 VGND VPWR sky130_fd_sc_hd__decap_12
X_5505_ _5501_/X _5502_/X _5503_/Y _5504_/X _5505_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_173_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_764 VGND VPWR sky130_fd_sc_hd__decap_8
X_6485_ _6426_/X _6484_/X _6481_/X _6485_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_3697_ wbs_we_i _3709_/C VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_134_937 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_1005 VGND VPWR sky130_fd_sc_hd__fill_2
X_5436_ _5372_/X _5373_/X _5372_/X _5373_/X _5436_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_134_959 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_5367_ _4461_/A _5123_/B _5367_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_87_501 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_288 VGND VPWR sky130_fd_sc_hd__decap_12
X_7106_ _7093_/X _7104_/X _7105_/Y _7631_/D VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_102_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_523 VGND VPWR sky130_fd_sc_hd__decap_12
X_4318_ _4200_/A _4200_/B _4200_/X _4318_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_141_480 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_171 VGND VPWR sky130_fd_sc_hd__decap_12
X_5298_ _5290_/X _5297_/X _5290_/X _5297_/X _5298_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7037_ _7037_/A _7037_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4249_ _4213_/X _4247_/X _4213_/X _4247_/X _4249_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_74_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1123 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_678 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_998 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_45 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_823 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_873 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_501 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_867 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_697 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1045 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_764 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_870 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_775 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1124 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_477 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_287 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_183_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_642 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_24_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_770 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1224 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_100 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1133 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_144 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_768 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_609 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_147 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_169 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_489 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1062 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1084 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_119_208 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1123 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_1027 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_881 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_560 VGND VPWR sky130_fd_sc_hd__decap_12
X_6270_ _5822_/X _5856_/B _5990_/X _6270_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_170_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1227 VGND VPWR sky130_fd_sc_hd__decap_12
X_5221_ _5089_/X _5090_/X _5089_/X _5090_/X _5221_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_103_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_1060 VGND VPWR sky130_fd_sc_hd__decap_8
X_5152_ _5136_/X _5151_/X _5136_/X _5151_/X _5152_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_29_1074 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_707 VGND VPWR sky130_fd_sc_hd__decap_12
X_4103_ _4098_/X _4099_/X _4102_/Y _4104_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_110_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_504 VGND VPWR sky130_fd_sc_hd__decap_12
X_5083_ _5078_/X _5082_/X _5078_/X _5082_/X _5083_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_1028 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_921 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_60 VGND VPWR sky130_fd_sc_hd__fill_1
X_4034_ _4032_/X _4034_/B _4035_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_38_965 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_93 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_762 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_732 VGND VPWR sky130_fd_sc_hd__decap_6
X_5985_ _5985_/A _5984_/Y _5985_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_109 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_428 VGND VPWR sky130_fd_sc_hd__decap_12
X_7724_ _6463_/X _6394_/A _7785_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_12_309 VGND VPWR sky130_fd_sc_hd__decap_12
X_4936_ _4868_/X _4869_/X _4850_/X _4870_/X _4936_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_40_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_642 VGND VPWR sky130_fd_sc_hd__decap_12
X_7655_ _6912_/X _6846_/A _7754_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA_10 _6219_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4867_ _4865_/X _4866_/X _4865_/X _4866_/X _4867_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_127_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_876 VGND VPWR sky130_fd_sc_hd__fill_2
X_6606_ _7694_/Q _6606_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_165_325 VGND VPWR sky130_fd_sc_hd__decap_12
X_3818_ _4646_/A _4547_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_7586_ _7586_/HI la_data_out[113] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_177_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_731 VGND VPWR sky130_fd_sc_hd__fill_1
X_4798_ _4540_/Y _4541_/X _4540_/Y _4541_/X _4798_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6537_ _6530_/A _6530_/B _6530_/X _6536_/X _6537_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_3749_ _5294_/A _3712_/X _3751_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_192_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_572 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_263 VGND VPWR sky130_fd_sc_hd__decap_12
X_6468_ _6466_/X _6468_/B _6467_/Y _6468_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_122_918 VGND VPWR sky130_fd_sc_hd__decap_12
X_5419_ _5360_/X _5364_/X _5360_/X _5364_/X _5419_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6399_ _6397_/Y _6398_/Y _6397_/Y _6398_/Y _6399_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_714 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1100 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_620 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_631 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_1193 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_865 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1087 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1038 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_898 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_1049 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_998 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_727 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_147 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1221 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_32 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_489 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_951 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_653 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_922 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_539 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_1189 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_825 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_292 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_346 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_520 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_1011 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_288 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_139_1099 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1244 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_334 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1054 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_464 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1034 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_497 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_294 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_417 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_179_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_776 VGND VPWR sky130_fd_sc_hd__decap_12
X_5770_ _5651_/X _5652_/X _5644_/X _5653_/X _5770_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_188_951 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_4721_ _4716_/X _4720_/X _4719_/X _4721_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_148_837 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_623 VGND VPWR sky130_fd_sc_hd__decap_6
X_7440_ io_oeb[35] _7440_/LO VGND VPWR sky130_fd_sc_hd__conb_1
X_4652_ _4645_/X _4651_/X _4645_/X _4651_/X _4652_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_159_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_645 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_859 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_818 VGND VPWR sky130_fd_sc_hd__decap_12
X_7371_ io_in[26] _7371_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_174_166 VGND VPWR sky130_fd_sc_hd__decap_12
X_4583_ _4583_/A _5533_/B _4583_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_116_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_317 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_626 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_572 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1081 VGND VPWR sky130_fd_sc_hd__decap_12
X_6322_ wbs_adr_i[1] wbs_adr_i[0] wbs_adr_i[3] _7258_/A _7264_/B VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_157_1111 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_391 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_5_0_wb_clk_i clkbuf_3_2_0_wb_clk_i/X _7756_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_196_1182 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_618 VGND VPWR sky130_fd_sc_hd__decap_12
X_6253_ _6240_/A _6253_/B _6253_/C _6255_/A VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_131_715 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1046 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1128 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_428 VGND VPWR sky130_fd_sc_hd__decap_12
X_5204_ _5137_/X _5141_/X _5137_/X _5141_/X _5204_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_170_394 VGND VPWR sky130_fd_sc_hd__decap_3
X_6184_ _6256_/B _6177_/X _6183_/Y _4888_/A _6073_/X _6185_/B VGND VPWR sky130_fd_sc_hd__o32a_4
X_5135_ _5133_/X _5134_/X _5133_/X _5134_/X _5135_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_111_461 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_995 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_835 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_537 VGND VPWR sky130_fd_sc_hd__decap_12
X_5066_ _5063_/X _5064_/X _5065_/X _5066_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_38_762 VGND VPWR sky130_fd_sc_hd__fill_1
X_4017_ _4625_/B _4748_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_42_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_389 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_935 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_1240 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_795 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1145 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1107 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1235 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_765 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_489 VGND VPWR sky130_fd_sc_hd__decap_8
X_5968_ _6319_/A _7730_/Q _7746_/Q _5968_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_201_708 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_973 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1123 VGND VPWR sky130_fd_sc_hd__decap_12
X_4919_ _4919_/A _4756_/B _4919_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7707_ _6576_/X _6507_/A _7707_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_40_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_601 VGND VPWR sky130_fd_sc_hd__decap_12
X_5899_ _5890_/X _5891_/X _5890_/X _5891_/X _5899_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_194_921 VGND VPWR sky130_fd_sc_hd__decap_12
X_7638_ _7022_/X _7638_/Q _7624_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_21_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_987 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_464 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_550 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_194 VGND VPWR sky130_fd_sc_hd__decap_12
X_7569_ _7569_/HI la_data_out[96] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_153_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_701 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_140_1170 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1154 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1048 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1176 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_1059 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_575 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_748 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_973 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_577 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_367 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_902 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_250 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_1245 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_726 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_1226 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_776 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_253 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_489 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_86 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_781 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_623 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_150 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1005 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_453 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_1240 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_604 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_380 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_851 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_152_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_726 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_459 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_1150 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1172 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_1055 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1036 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1058 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_507 VGND VPWR sky130_fd_sc_hd__decap_12
X_6940_ _6940_/A _6940_/B _6940_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_82_849 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_874 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_294 VGND VPWR sky130_fd_sc_hd__decap_8
X_6871_ _6840_/Y _6842_/B _6842_/X _6870_/X _6871_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_23_916 VGND VPWR sky130_fd_sc_hd__fill_2
X_5822_ _5815_/X _5816_/X _5815_/X _5816_/X _5822_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_23_927 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_269 VGND VPWR sky130_fd_sc_hd__decap_12
X_5753_ _5749_/X _5750_/X _5751_/Y _5752_/X _5753_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_22_459 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_921 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1173 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1004 VGND VPWR sky130_fd_sc_hd__decap_12
X_4704_ _4558_/X _4559_/X _4558_/X _4559_/X _4704_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_194_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1195 VGND VPWR sky130_fd_sc_hd__decap_12
X_5684_ _5684_/A _5684_/B _5684_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_136_807 VGND VPWR sky130_fd_sc_hd__decap_12
X_7423_ io_oeb[18] _7423_/LO VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_148_678 VGND VPWR sky130_fd_sc_hd__decap_12
X_4635_ _4634_/A _4634_/B _4634_/X _4635_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_135_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1119 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_7354_ _7354_/A _7354_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_128_380 VGND VPWR sky130_fd_sc_hd__decap_12
X_4566_ _4566_/A _4565_/X _4581_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_2_809 VGND VPWR sky130_fd_sc_hd__decap_12
X_6305_ _6299_/Y _6300_/Y _6305_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_144_873 VGND VPWR sky130_fd_sc_hd__decap_12
X_7285_ _7749_/Q _7280_/X _7281_/X _7284_/Y wbs_dat_o[3] VGND VPWR sky130_fd_sc_hd__a211o_4
X_4497_ _5304_/A _4497_/B _4497_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_104_726 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_523 VGND VPWR sky130_fd_sc_hd__decap_12
X_6236_ _6308_/B _6240_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_134_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1160 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_269 VGND VPWR sky130_fd_sc_hd__fill_1
X_6167_ _6165_/Y _6166_/X _6167_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_135_1261 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_621 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_1166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_1008 VGND VPWR sky130_fd_sc_hd__decap_12
X_5118_ _5091_/X _5106_/X _5116_/X _5117_/X _5118_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_58_868 VGND VPWR sky130_fd_sc_hd__decap_12
X_6098_ _6097_/X _6098_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_100_987 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_367 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_35 VGND VPWR sky130_fd_sc_hd__decap_12
X_5049_ _5042_/X _5048_/X _5050_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_73_838 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_710 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_337 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_754 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_220 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_534 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_415 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_297 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_45 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_971 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1224 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1268 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_998 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_810 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1093 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_831 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_854 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_1047 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_864 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1244 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_602 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_676 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_581 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_1031 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_1046 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_668 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_1068 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_724 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1097 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_1067 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_910 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_245 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_270 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_239 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_281 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_292 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_964 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_604 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_829 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_475 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_423 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_957 VGND VPWR sky130_fd_sc_hd__decap_12
X_4420_ _4418_/X _4419_/X _4418_/X _4419_/X _4420_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1111 VGND VPWR sky130_fd_sc_hd__decap_12
X_4351_ _4347_/X _4350_/X _4347_/X _4350_/X _4351_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_724 VGND VPWR sky130_fd_sc_hd__decap_8
X_7070_ _7070_/A _7070_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4282_ _4280_/X _4281_/X _4279_/X _4282_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_193_1196 VGND VPWR sky130_fd_sc_hd__decap_12
X_6021_ _5050_/A _6020_/Y _6021_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_113_578 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_952 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_985 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_495 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1240 VGND VPWR sky130_fd_sc_hd__decap_8
X_6923_ _6923_/A _6862_/X _6923_/C _7651_/D VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_78_1262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6854_ _6852_/Y _6853_/Y _6854_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_126_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_234 VGND VPWR sky130_fd_sc_hd__decap_8
X_5805_ _5794_/X _5805_/B _5805_/X VGND VPWR sky130_fd_sc_hd__and2_4
XPHY_1808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6785_ _6670_/A _6785_/X VGND VPWR sky130_fd_sc_hd__buf_1
XPHY_1819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3997_ _3997_/A _4027_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_195_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_565 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_869 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_5736_ _4697_/A _4482_/A _5736_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_129_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_475 VGND VPWR sky130_fd_sc_hd__decap_12
X_5667_ _5590_/X _5597_/B _5597_/X _5667_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_129_59 VGND VPWR sky130_fd_sc_hd__fill_2
X_4618_ _4568_/X _4572_/X _4571_/X _4618_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_7406_ io_oeb[1] _7406_/LO VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_50_1181 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_1036 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_1143 VGND VPWR sky130_fd_sc_hd__decap_12
X_5598_ _4455_/A _4778_/B _5598_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_135_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_851 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_70 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_607 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_618 VGND VPWR sky130_fd_sc_hd__decap_12
X_7337_ _5632_/A _7309_/X _7332_/X _7336_/Y wbs_dat_o[12] VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_163_489 VGND VPWR sky130_fd_sc_hd__decap_8
X_4549_ _4549_/A _4549_/B _4549_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_104_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_681 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_821 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_1203 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_692 VGND VPWR sky130_fd_sc_hd__decap_8
X_7268_ _7746_/Q _7257_/X _7260_/X _7267_/Y wbs_dat_o[0] VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_89_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_919 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_353 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_407 VGND VPWR sky130_fd_sc_hd__decap_12
X_6219_ _6219_/A _6219_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_132_898 VGND VPWR sky130_fd_sc_hd__decap_12
X_7199_ _7154_/Y _7155_/Y _7156_/X _7198_/X _7199_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_86_963 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_56 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_67 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_153 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_484 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_1250 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_646 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_337 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_810 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_178 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_746 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_245 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_289 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1160 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_773 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1073 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_1024 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_935 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1046 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_1136 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_681 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_407 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_386 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_1172 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1025 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1119 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_698 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_337 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1118 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_540 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_999 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_487 VGND VPWR sky130_fd_sc_hd__fill_1
X_3920_ _4648_/A _4743_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_51_329 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_696 VGND VPWR sky130_fd_sc_hd__decap_12
X_3851_ _3850_/Y _4680_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_6570_ _6549_/X _6568_/X _6569_/Y _7709_/D VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_81_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_3782_ wbs_dat_i[15] _3790_/B _3782_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_34_1154 VGND VPWR sky130_fd_sc_hd__decap_4
X_5521_ _4800_/X _4801_/X _4800_/X _4801_/X _5521_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_9_761 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_795 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_1184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_1135 VGND VPWR sky130_fd_sc_hd__decap_12
X_5452_ _5400_/X _5440_/X _5450_/X _5451_/X _5452_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_117_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_916 VGND VPWR sky130_fd_sc_hd__decap_12
X_4403_ _4401_/X _4402_/X _4401_/X _4402_/X _4403_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_195_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_489 VGND VPWR sky130_fd_sc_hd__decap_3
X_5383_ _5383_/A _5383_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_132_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_821 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_532 VGND VPWR sky130_fd_sc_hd__decap_12
X_7122_ _7085_/X _7121_/X _7114_/X _7122_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_119_1020 VGND VPWR sky130_fd_sc_hd__decap_12
X_4334_ _4844_/A _4591_/B _4336_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_160_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_640 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_865 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_554 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1008 VGND VPWR sky130_fd_sc_hd__decap_8
X_7053_ la_data_in[88] _7053_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_141_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_898 VGND VPWR sky130_fd_sc_hd__decap_12
X_4265_ _4264_/A _4263_/X _4264_/X _4265_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_99_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1130 VGND VPWR sky130_fd_sc_hd__fill_1
X_6004_ _5566_/X _6004_/B _6004_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_41_1103 VGND VPWR sky130_fd_sc_hd__fill_1
X_4196_ _4156_/X _4193_/X _4194_/X _4195_/X _4196_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_83_900 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_602 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_175 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_966 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_605 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_871 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_178 VGND VPWR sky130_fd_sc_hd__decap_4
X_6906_ _6870_/X _6904_/X _6905_/X _6906_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_42_329 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_830 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_863 VGND VPWR sky130_fd_sc_hd__decap_3
X_6837_ _6837_/A _6837_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_1605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_633 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_215 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_154 VGND VPWR sky130_fd_sc_hd__decap_12
X_6768_ _6717_/A _6717_/B _6717_/X _6767_/X _6768_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_10_226 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1081 VGND VPWR sky130_fd_sc_hd__decap_12
X_5719_ _5678_/X _5717_/X _5678_/X _5717_/X _5719_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6699_ _6633_/A la_data_in[19] _6635_/X _6699_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_176_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_423 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_968 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_562 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_404 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_960 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1085 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_727 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_900 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_944 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_207_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_281 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_443 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1152 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_999 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_98 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_318 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1105 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_543 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_515 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_684 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1045 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_633 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_340 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1067 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1089 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_86 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_489 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_681 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1100 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_993 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_824 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_695 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_546 VGND VPWR sky130_fd_sc_hd__decap_12
X_4050_ _3722_/A _4925_/B _4050_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_49_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_900 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_378 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1051 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_145 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_307 VGND VPWR sky130_fd_sc_hd__decap_8
X_4952_ _4951_/X _4952_/B _4952_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7740_ _6347_/Y _7740_/Q _7806_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_75_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_498 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_983 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_392 VGND VPWR sky130_fd_sc_hd__decap_12
X_3903_ _5200_/A _5215_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_51_159 VGND VPWR sky130_fd_sc_hd__decap_12
X_4883_ _4881_/Y _4883_/B _4883_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_7671_ _7671_/D _7671_/Q _7756_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_36_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_334 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_682 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_373 VGND VPWR sky130_fd_sc_hd__decap_12
X_3834_ _4656_/A _4455_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_6622_ la_data_in[23] _6623_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_177_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1221 VGND VPWR sky130_fd_sc_hd__decap_12
X_6553_ _6560_/A _6553_/B _6553_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_146_710 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_568 VGND VPWR sky130_fd_sc_hd__decap_12
X_3765_ _4498_/A _4503_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_158_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1090 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_423 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_220 VGND VPWR sky130_fd_sc_hd__decap_12
X_5504_ _5501_/X _5502_/X _5501_/X _5502_/X _5504_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_754 VGND VPWR sky130_fd_sc_hd__decap_8
X_6484_ _7716_/Q la_data_in[114] _6420_/X _6484_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_3696_ wbs_cyc_i wbs_stb_i _6038_/B VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_106_607 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_562 VGND VPWR sky130_fd_sc_hd__decap_12
X_5435_ _5413_/X _5414_/X _5407_/X _5415_/X _5435_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_161_724 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_195_1099 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_1203 VGND VPWR sky130_fd_sc_hd__decap_6
X_5366_ _4645_/A _4778_/B _5366_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_142_971 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_204 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_929 VGND VPWR sky130_fd_sc_hd__fill_1
X_4317_ _4316_/A _4315_/X _4447_/B _4317_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_7105_ _7093_/X _7104_/X _7024_/X _7105_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_82_1258 VGND VPWR sky130_fd_sc_hd__fill_1
X_5297_ _5291_/X _5296_/X _5291_/X _5296_/X _5297_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_87_535 VGND VPWR sky130_fd_sc_hd__decap_12
X_7036_ _7034_/Y _7035_/Y _7034_/Y _7035_/Y _7095_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_4248_ _7779_/Q _4248_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_206_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_101 VGND VPWR sky130_fd_sc_hd__decap_12
X_4179_ _4179_/A _4179_/B _4179_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_67_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_808 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_413 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_318 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_958 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_690 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_446 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1143 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_835 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_513 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_345 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_654 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_208_1187 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_507 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_401 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_849 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_754 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_540 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1057 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1079 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_882 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_787 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_178_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1109 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_448 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_459 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_245 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_684 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_676 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1161 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1236 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_112 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1145 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1205 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_966 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_1028 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1118 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_487 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_947 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_4050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_964 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1096 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_192 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1162 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_337 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1252 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_702 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_893 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_572 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_532 VGND VPWR sky130_fd_sc_hd__decap_12
X_5220_ _5214_/X _5217_/X _5218_/X _5219_/X _5220_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_192_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_971 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1114 VGND VPWR sky130_fd_sc_hd__fill_1
X_5151_ _5142_/X _5148_/X _5149_/X _5150_/X _5151_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_96_310 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1086 VGND VPWR sky130_fd_sc_hd__decap_12
X_4102_ _4102_/A _4102_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_9_1169 VGND VPWR sky130_fd_sc_hd__decap_8
X_5082_ _5079_/X _5080_/X _5081_/X _5082_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_57_719 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1067 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1018 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_516 VGND VPWR sky130_fd_sc_hd__decap_3
X_4033_ _3991_/A _3990_/X _3991_/X _4034_/B VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_96_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_933 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_741 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_785 VGND VPWR sky130_fd_sc_hd__decap_8
X_5984_ _5941_/X _5942_/X _5983_/X _5984_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_52_457 VGND VPWR sky130_fd_sc_hd__fill_1
X_7723_ _7723_/D _7723_/Q _7785_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_468 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1002 VGND VPWR sky130_fd_sc_hd__decap_4
X_4935_ _4922_/X _4934_/X _4922_/X _4934_/X _4935_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_162_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_654 VGND VPWR sky130_fd_sc_hd__decap_12
X_7654_ _7654_/D _7654_/Q _7754_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA_11 _6319_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_4866_ _4645_/X _4651_/X _4650_/X _4866_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_127_1196 VGND VPWR sky130_fd_sc_hd__decap_12
X_6605_ _6605_/A _6605_/B _6605_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_123_1038 VGND VPWR sky130_fd_sc_hd__decap_12
X_3817_ _7804_/Q _4646_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_193_635 VGND VPWR sky130_fd_sc_hd__decap_12
X_4797_ _4786_/X _4787_/X _4785_/X _4788_/X _4797_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_7585_ _7585_/HI la_data_out[112] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_165_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1062 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_398 VGND VPWR sky130_fd_sc_hd__decap_6
X_3748_ _4568_/A _5294_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_6536_ _6531_/Y _6532_/Y _6535_/X _6536_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_137_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_178 VGND VPWR sky130_fd_sc_hd__decap_12
X_6467_ _6467_/A _6467_/B _6467_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_137_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_448 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_459 VGND VPWR sky130_fd_sc_hd__decap_6
X_5418_ _5416_/X _5417_/X _5418_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_6398_ la_data_in[121] _6398_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_88_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_726 VGND VPWR sky130_fd_sc_hd__decap_12
X_5349_ _5157_/A _4757_/B _5349_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_134_1112 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1044 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1172 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_877 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_985 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1000 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1178 VGND VPWR sky130_fd_sc_hd__decap_12
X_7019_ _6955_/X _7019_/B _7019_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_29_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_914 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_739 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_159 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1113 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_800 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_44 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_963 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_665 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_934 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_804 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_343 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_624 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_837 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_495 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_337 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_336 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_172_808 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_510 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_757 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_971 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_855 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1248 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_719 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_398 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_538 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_590 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_346 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1044 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1066 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_560 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_251 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_424 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1005 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_1016 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_788 VGND VPWR sky130_fd_sc_hd__decap_12
X_4720_ _4717_/X _4718_/X _4719_/X _4720_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_187_440 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_3190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_602 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_816 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_794 VGND VPWR sky130_fd_sc_hd__decap_12
X_4651_ _4647_/X _4649_/X _4650_/X _4651_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_175_657 VGND VPWR sky130_fd_sc_hd__decap_12
X_4582_ _5294_/B _5533_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_7370_ _7370_/A _7370_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_190_605 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_329 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_190_638 VGND VPWR sky130_fd_sc_hd__decap_3
X_6321_ wbs_adr_i[2] _7258_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_122_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_391 VGND VPWR sky130_fd_sc_hd__decap_6
X_6252_ _6246_/Y _6250_/X _6253_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_115_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_362 VGND VPWR sky130_fd_sc_hd__decap_12
X_5203_ _5198_/X _5202_/X _5201_/X _5203_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_192_1058 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_6183_ _6174_/Y _6176_/X _6183_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_5134_ _5093_/X _5097_/X _5096_/X _5134_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_85_847 VGND VPWR sky130_fd_sc_hd__decap_6
X_5065_ _5063_/X _5064_/X _5065_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_123_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_869 VGND VPWR sky130_fd_sc_hd__decap_8
X_4016_ _4016_/A _4625_/B VGND VPWR sky130_fd_sc_hd__buf_1
XPHY_4808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_880 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_947 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_168_1252 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_1214 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_969 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_727 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1119 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_1247 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_777 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_928 VGND VPWR sky130_fd_sc_hd__decap_3
X_5967_ _7747_/Q _5966_/X _5958_/X _5967_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_52_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_980 VGND VPWR sky130_fd_sc_hd__decap_6
X_7706_ _6578_/X _6510_/A _7696_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4918_ _4915_/X _4916_/X _4917_/X _4918_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_179_985 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_205_1135 VGND VPWR sky130_fd_sc_hd__decap_12
X_5898_ _3901_/X _4363_/A _5898_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_166_613 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_933 VGND VPWR sky130_fd_sc_hd__decap_12
X_7637_ _7026_/X _7637_/Q _7624_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4849_ _4840_/X _4848_/X _4840_/X _4848_/X _4849_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_165_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_696 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_860 VGND VPWR sky130_fd_sc_hd__decap_12
X_7568_ _7568_/HI la_data_out[95] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_194_999 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_818 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_713 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1182 VGND VPWR sky130_fd_sc_hd__decap_8
X_6519_ _7703_/Q _6519_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_88_1264 VGND VPWR sky130_fd_sc_hd__decap_12
X_7499_ _7499_/HI la_data_out[26] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_134_532 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_107_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1128 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_771 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_825 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_996 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1150 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_828 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_560 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_711 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_402 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_265 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1249 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_98 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_98 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_602 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_410 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1044 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_162 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_111 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_977 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_184 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_616 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_678 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_587 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1050 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_685 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1067 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_886 VGND VPWR sky130_fd_sc_hd__decap_6
X_6870_ _6843_/Y _6844_/Y _6845_/X _6869_/X _6870_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_50_703 VGND VPWR sky130_fd_sc_hd__decap_12
X_5821_ _5821_/A _6269_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_23_939 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_980 VGND VPWR sky130_fd_sc_hd__decap_12
X_5752_ _5749_/X _5750_/X _5749_/X _5750_/X _5752_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_188_760 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1065 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_1016 VGND VPWR sky130_fd_sc_hd__decap_12
X_4703_ _4694_/X _4700_/X _4701_/X _4702_/X _4703_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_187_281 VGND VPWR sky130_fd_sc_hd__decap_12
X_5683_ _3877_/A _4901_/A _5684_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_176_955 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1008 VGND VPWR sky130_fd_sc_hd__decap_3
X_7422_ io_oeb[17] _7422_/LO VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_136_819 VGND VPWR sky130_fd_sc_hd__decap_4
X_4634_ _4634_/A _4634_/B _4634_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_135_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_649 VGND VPWR sky130_fd_sc_hd__decap_12
X_4565_ _4565_/A _4565_/B _4565_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7353_ _5383_/A _7388_/A _7348_/X _7352_/Y wbs_dat_o[15] VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_190_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_392 VGND VPWR sky130_fd_sc_hd__decap_4
X_6304_ _6211_/A _6304_/B _7750_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_116_554 VGND VPWR sky130_fd_sc_hd__decap_12
X_4496_ _4495_/A _4495_/B _4495_/X _4496_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_7284_ _5185_/A _7262_/X _7283_/X _7284_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_1_309 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_738 VGND VPWR sky130_fd_sc_hd__decap_12
X_6235_ _6211_/A _6234_/Y _7764_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_131_535 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_6166_ _5048_/X _6152_/X _5046_/X _6166_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_85_611 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_825 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_1273 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_922 VGND VPWR sky130_fd_sc_hd__decap_12
X_5117_ _5091_/X _5106_/X _5091_/X _5106_/X _5117_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_69_184 VGND VPWR sky130_fd_sc_hd__decap_12
X_6097_ _4210_/X _6096_/X _4205_/B _6097_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_44_1189 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_806 VGND VPWR sky130_fd_sc_hd__fill_1
X_5048_ _5045_/A _5045_/B _5047_/Y _5048_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_84_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1172 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_316 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_47 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_593 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_349 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_232 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1093 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_546 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1272 VGND VPWR sky130_fd_sc_hd__decap_4
X_6999_ _6905_/A _6999_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_40_224 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_900 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1236 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_983 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1258 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_977 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1001 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_852 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_18 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_682 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1067 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1059 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_342 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_876 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1207 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_397 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_292 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_666 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_806 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_688 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1036 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_861 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_574 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_894 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_950 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_260 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_257 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_271 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_282 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_421 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_281 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_293 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_741 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_999 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_785 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_1060 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_969 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_32_1093 VGND VPWR sky130_fd_sc_hd__decap_6
X_4350_ _4348_/X _4349_/X _4348_/X _4349_/X _4350_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_67_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_660 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1118 VGND VPWR sky130_fd_sc_hd__decap_8
X_4281_ _3722_/A _4459_/B _4281_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_101_708 VGND VPWR sky130_fd_sc_hd__decap_12
X_6020_ _5041_/X _5047_/Y _6019_/X _6020_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_79_460 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_611 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_140_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_379 VGND VPWR sky130_fd_sc_hd__decap_12
X_6922_ _6922_/A _6861_/X _6923_/C VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_54_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_530 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1252 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1274 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1233 VGND VPWR sky130_fd_sc_hd__decap_12
X_6853_ la_data_in[51] _6853_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_63_883 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_371 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1138 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_596 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_213 VGND VPWR sky130_fd_sc_hd__fill_1
X_5804_ _5727_/X _5746_/X _5747_/X _5804_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_161_1108 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1239 VGND VPWR sky130_fd_sc_hd__decap_12
X_6784_ _6718_/A la_data_in[43] _6720_/X _6784_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_23_769 VGND VPWR sky130_fd_sc_hd__decap_12
X_3996_ _3988_/Y _3989_/X _3988_/Y _3989_/X _3996_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_50_577 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_410 VGND VPWR sky130_fd_sc_hd__decap_12
X_5735_ _5730_/X _5734_/X _5733_/X _5735_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_22_279 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1116 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_977 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_988 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_27 VGND VPWR sky130_fd_sc_hd__decap_12
X_5666_ _3904_/X _4126_/B _5668_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_148_487 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1111 VGND VPWR sky130_fd_sc_hd__decap_3
X_7405_ io_oeb[0] _7405_/LO VGND VPWR sky130_fd_sc_hd__conb_1
X_4617_ _4612_/X _4616_/X _4612_/X _4616_/X _4617_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_117_830 VGND VPWR sky130_fd_sc_hd__fill_2
X_5597_ _5590_/X _5597_/B _5597_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_209_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1155 VGND VPWR sky130_fd_sc_hd__decap_4
X_7336_ _4589_/A _7322_/X _7335_/X _7336_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
X_4548_ _4548_/A _4591_/B _4549_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_172_980 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_513 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_150_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_7267_ _3904_/X _7262_/X _7266_/X _7267_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_145_59 VGND VPWR sky130_fd_sc_hd__fill_2
X_4479_ _4479_/A _4479_/B _4486_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_89_257 VGND VPWR sky130_fd_sc_hd__decap_12
X_6218_ _6214_/Y _6215_/X _6217_/X _6218_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_131_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_419 VGND VPWR sky130_fd_sc_hd__decap_8
X_7198_ _7157_/Y _7158_/Y _7225_/B _7198_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_131_387 VGND VPWR sky130_fd_sc_hd__fill_1
X_6149_ _4807_/X _6149_/B _6150_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_100_741 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_752 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_79 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_165 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_891 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_4413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1008 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_349 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_861 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_703 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_522 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_758 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_190 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_217 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_741 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1044 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1036 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1058 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1148 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_693 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_150_630 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_706 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_888 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_419 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1151 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_964 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_458 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_1244 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_469 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1138 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_135 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_669 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_544 VGND VPWR sky130_fd_sc_hd__decap_12
X_3850_ _3850_/A _3850_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_73_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_886 VGND VPWR sky130_fd_sc_hd__decap_12
X_3781_ _4552_/A _3767_/B _3781_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_160_1130 VGND VPWR sky130_fd_sc_hd__decap_12
X_5520_ _6198_/A _6198_/B _6000_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_201_881 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_402 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_773 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_273 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_733 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_744 VGND VPWR sky130_fd_sc_hd__decap_12
X_5451_ _5400_/X _5440_/X _5400_/X _5440_/X _5451_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_201_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_159 VGND VPWR sky130_fd_sc_hd__decap_12
X_4402_ _5058_/A _4923_/B _4402_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_161_928 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_939 VGND VPWR sky130_fd_sc_hd__decap_12
X_5382_ _4552_/A _4793_/B _5382_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_172_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_511 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_7121_ _7055_/A la_data_in[87] _7057_/X _7121_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_4333_ _4328_/X _4332_/X _4331_/X _4333_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_119_1032 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_652 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1054 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_877 VGND VPWR sky130_fd_sc_hd__decap_8
X_4264_ _4264_/A _4263_/X _4264_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7052_ _7626_/Q _7052_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_113_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_588 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_141_696 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_227 VGND VPWR sky130_fd_sc_hd__decap_12
X_6003_ _5575_/X _5581_/Y _6002_/X _6004_/B VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_39_110 VGND VPWR sky130_fd_sc_hd__decap_12
X_4195_ _4187_/X _4190_/Y _4186_/X _4191_/X _4195_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_68_986 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_485 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_992 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_989 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_617 VGND VPWR sky130_fd_sc_hd__decap_12
X_6905_ _6905_/A _6905_/X VGND VPWR sky130_fd_sc_hd__buf_1
XPHY_3019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1060 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_883 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_803 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_393 VGND VPWR sky130_fd_sc_hd__decap_8
X_6836_ _6834_/Y _6835_/Y _6834_/Y _6835_/Y _6874_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_2329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1014 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1066 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_94 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_645 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_869 VGND VPWR sky130_fd_sc_hd__decap_12
X_6767_ _6720_/A _6720_/B _6720_/X _6766_/X _6767_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XPHY_1639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1069 VGND VPWR sky130_fd_sc_hd__decap_12
X_3979_ _3972_/X _3979_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_50_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_238 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_379 VGND VPWR sky130_fd_sc_hd__decap_12
X_5718_ _5712_/X _5713_/X _5711_/Y _5714_/X _5718_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_206_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_251 VGND VPWR sky130_fd_sc_hd__decap_12
X_6698_ _6694_/X _6698_/B _6697_/Y _7686_/D VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_176_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_435 VGND VPWR sky130_fd_sc_hd__decap_4
X_5649_ _5605_/X _5611_/X _5604_/X _5612_/X _5649_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_163_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_541 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_799 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_416 VGND VPWR sky130_fd_sc_hd__decap_8
X_7319_ _5751_/A _7309_/X _7315_/X _7318_/Y wbs_dat_o[9] VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_85_1053 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_855 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_459 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1097 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1067 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_912 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_986 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_496 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_113 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_809 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_455 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1142 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_105 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1141 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_555 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1174 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1245 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_352 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_886 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_98 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_906 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_794 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_671 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_693 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1134 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_814 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_836 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_558 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_912 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_794 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_135 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_1063 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_617 VGND VPWR sky130_fd_sc_hd__decap_12
X_4951_ _4947_/X _4950_/Y _4947_/X _4950_/Y _4951_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_75_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_995 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_842 VGND VPWR sky130_fd_sc_hd__decap_12
X_3902_ _3901_/X _5200_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_162_1203 VGND VPWR sky130_fd_sc_hd__decap_8
X_7670_ _6805_/X _7670_/Q _7756_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_178_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_190 VGND VPWR sky130_fd_sc_hd__decap_12
X_4882_ _4880_/X _4883_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_177_324 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1239 VGND VPWR sky130_fd_sc_hd__decap_12
X_6621_ _7689_/Q _6621_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_3833_ _7802_/Q _4656_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_177_346 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_379 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_1233 VGND VPWR sky130_fd_sc_hd__decap_12
X_6552_ _6495_/Y _6496_/Y _6497_/X _6551_/X _6553_/B VGND VPWR sky130_fd_sc_hd__o22a_4
X_3764_ _4570_/A _4498_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_158_593 VGND VPWR sky130_fd_sc_hd__decap_4
X_5503_ _5503_/A _5503_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_192_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_435 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1001 VGND VPWR sky130_fd_sc_hd__decap_12
X_6483_ _6427_/X _6479_/X _6482_/Y _7717_/D VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_145_232 VGND VPWR sky130_fd_sc_hd__decap_12
X_3695_ _3695_/A _6038_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_12_1250 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_405 VGND VPWR sky130_fd_sc_hd__decap_12
X_5434_ _5419_/X _5425_/X _5432_/X _5433_/X _5434_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_173_574 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_330 VGND VPWR sky130_fd_sc_hd__decap_12
X_5365_ _5360_/X _5364_/X _5363_/X _5365_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_102_803 VGND VPWR sky130_fd_sc_hd__decap_12
X_7104_ _7037_/A la_data_in[93] _7039_/X _7104_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_4316_ _4316_/A _4315_/X _4447_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_142_983 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_216 VGND VPWR sky130_fd_sc_hd__decap_12
X_5296_ _5292_/Y _5295_/X _5292_/Y _5295_/X _5296_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_102_836 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_847 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_7035_ la_data_in[94] _7035_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4247_ _4214_/X _4244_/X _4245_/X _4246_/X _4247_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_68_761 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_142_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1040 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_379 VGND VPWR sky130_fd_sc_hd__decap_12
X_4178_ _4565_/A _4235_/B _4179_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_56_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_113 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_1158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_948 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_639 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_425 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_814 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_0_0_wb_clk_i clkbuf_1_0_1_wb_clk_i/X clkbuf_2_0_1_wb_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_2115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1155 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_352 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_847 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_633 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_886 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_672 VGND VPWR sky130_fd_sc_hd__decap_12
X_6819_ _6819_/A _6819_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_525 VGND VPWR sky130_fd_sc_hd__decap_12
X_7799_ _7799_/D _3858_/A _7801_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1199 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_1030 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_497 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_518 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_413 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1036 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1039 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_201 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_757 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_3 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_768 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_279 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_471 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_208 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_688 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1211 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_794 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_411 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1173 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1248 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_124 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_737 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_1157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1217 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_1228 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_989 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_4040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_93 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1258 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_425 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_4062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_853 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_611 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_80 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_661 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_91 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_823 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_806 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_396 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_828 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1231 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_733 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_349 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_744 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_714 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_788 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_980 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1010 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_983 VGND VPWR sky130_fd_sc_hd__decap_12
X_5150_ _5142_/X _5148_/X _5142_/X _5148_/X _5150_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_116_1002 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_780 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_633 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_322 VGND VPWR sky130_fd_sc_hd__decap_12
X_4101_ _4101_/A _4102_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_155_1084 VGND VPWR sky130_fd_sc_hd__decap_12
X_5081_ _5079_/X _5080_/X _5081_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_97_867 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_154 VGND VPWR sky130_fd_sc_hd__decap_12
X_4032_ _3996_/X _4031_/X _4032_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_111_688 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_84 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_444 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_550 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_105 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_425 VGND VPWR sky130_fd_sc_hd__decap_12
X_5983_ _5983_/A _6293_/B _5983_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_24_138 VGND VPWR sky130_fd_sc_hd__decap_12
X_7722_ _6468_/X _6400_/A _7785_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4934_ _4932_/X _4933_/X _4932_/X _4933_/X _4934_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_166_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_672 VGND VPWR sky130_fd_sc_hd__decap_12
X_7653_ _6918_/X _7653_/Q _7756_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_162_1044 VGND VPWR sky130_fd_sc_hd__decap_12
X_4865_ _4860_/X _4864_/X _4860_/X _4864_/X _4865_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_178_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_491 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_12 _6319_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_1069 VGND VPWR sky130_fd_sc_hd__decap_12
X_6604_ la_data_in[29] _6605_/B VGND VPWR sky130_fd_sc_hd__inv_8
X_3816_ _3791_/A _3814_/X _3815_/Y _3816_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_7584_ _7584_/HI la_data_out[111] VGND VPWR sky130_fd_sc_hd__conb_1
X_4796_ _4792_/X _4793_/X _4794_/Y _4795_/X _4796_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_159_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_388 VGND VPWR sky130_fd_sc_hd__decap_8
X_6535_ _6596_/A _6596_/B _6535_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_3747_ _4919_/A _4568_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_203_1074 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_703 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_928 VGND VPWR sky130_fd_sc_hd__decap_8
X_6466_ _6595_/A _6466_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_174_894 VGND VPWR sky130_fd_sc_hd__fill_1
X_5417_ _5339_/X _5345_/X _5346_/X _5417_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_6397_ _7723_/Q _6397_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_133_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1170 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_705 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_419 VGND VPWR sky130_fd_sc_hd__decap_8
X_5348_ _5348_/A _4758_/B _5348_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_114_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_738 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_1124 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_749 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_655 VGND VPWR sky130_fd_sc_hd__decap_12
X_5279_ _5274_/X _5276_/X _5277_/Y _5278_/X _5279_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_153_59 VGND VPWR sky130_fd_sc_hd__fill_2
X_7018_ _6976_/X _7016_/X _7017_/Y _7640_/D VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_130_997 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_1012 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1209 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_904 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_989 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_712 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_926 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_909 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_425 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_611 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_812 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_56 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_975 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_261 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_816 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_355 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_636 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_849 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_135 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_703 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_714 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_265 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_510 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1210 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_886 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_823 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_344 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_709 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_485 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_1180 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_572 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_414 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_436 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_672 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_642 VGND VPWR sky130_fd_sc_hd__decap_8
X_4650_ _4647_/X _4649_/X _4650_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_2490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_496 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_669 VGND VPWR sky130_fd_sc_hd__fill_2
X_4581_ _4581_/A _4581_/B _4581_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_6320_ _6332_/A _6320_/B _6319_/X _7746_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_171_853 VGND VPWR sky130_fd_sc_hd__fill_1
X_6251_ _6246_/Y _6250_/X _6253_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_182_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_257 VGND VPWR sky130_fd_sc_hd__decap_4
X_5202_ _5199_/X _5201_/B _5201_/X _5202_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_170_374 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_588 VGND VPWR sky130_fd_sc_hd__decap_12
X_6182_ _6179_/X _6180_/Y _6181_/X _7773_/D VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_124_780 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_227 VGND VPWR sky130_fd_sc_hd__decap_12
X_5133_ _5128_/X _5132_/X _5128_/X _5132_/X _5133_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_141 VGND VPWR sky130_fd_sc_hd__decap_12
X_5064_ _4553_/A _4485_/B _5064_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_42_1040 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_496 VGND VPWR sky130_fd_sc_hd__decap_12
X_4015_ _7741_/Q _4016_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_65_550 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_520 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_391 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_745 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_164_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_739 VGND VPWR sky130_fd_sc_hd__decap_12
X_5966_ _7795_/Q _7730_/Q _5966_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_53_789 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_1261 VGND VPWR sky130_fd_sc_hd__decap_3
X_7705_ _6581_/X _7705_/Q _7696_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_288 VGND VPWR sky130_fd_sc_hd__decap_12
X_4917_ _4915_/X _4916_/X _4917_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_139_806 VGND VPWR sky130_fd_sc_hd__decap_12
X_5897_ _5870_/X _5871_/X _5872_/X _5897_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_32_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_305 VGND VPWR sky130_fd_sc_hd__decap_12
X_7636_ _7029_/X _7636_/Q _7624_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_166_625 VGND VPWR sky130_fd_sc_hd__decap_12
X_4848_ _4846_/X _4847_/X _4846_/X _4847_/X _4848_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_20_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1142 VGND VPWR sky130_fd_sc_hd__decap_12
X_7567_ _7567_/HI la_data_out[94] VGND VPWR sky130_fd_sc_hd__conb_1
X_4779_ _4779_/A _4779_/B _4779_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_147_872 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_6518_ _6516_/Y _6518_/B _6518_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_107_725 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_318 VGND VPWR sky130_fd_sc_hd__decap_12
X_7498_ _7498_/HI la_data_out[25] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_88_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_769 VGND VPWR sky130_fd_sc_hd__decap_12
X_6449_ _6449_/A _6442_/X _6450_/C VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_122_706 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_363 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_441 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_804 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_557 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_783 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_314 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_309 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_336 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1162 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_807 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_572 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1168 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_1206 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_918 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_277 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_420 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_428 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_620 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1001 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_642 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_794 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_984 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_809 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_174 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_123 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_989 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_861 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_511 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_831 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_697 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_794 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1106 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_678 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_550 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_274 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_745 VGND VPWR sky130_fd_sc_hd__decap_12
X_5820_ _5820_/A _5819_/X _5821_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_50_715 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_992 VGND VPWR sky130_fd_sc_hd__decap_12
X_5751_ _5751_/A _5751_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_210_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_1191 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_951 VGND VPWR sky130_fd_sc_hd__decap_8
X_4702_ _4694_/X _4700_/X _4694_/X _4700_/X _4702_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_203_581 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_934 VGND VPWR sky130_fd_sc_hd__decap_12
X_5682_ _5178_/A _4291_/A _5684_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_33_1028 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_293 VGND VPWR sky130_fd_sc_hd__decap_12
X_7421_ io_oeb[16] _7421_/LO VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_147_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_483 VGND VPWR sky130_fd_sc_hd__decap_4
X_4633_ _3778_/A _4145_/A _4634_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_124_1189 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1219 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_7352_ _4552_/A _7349_/X _7351_/X _7352_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_200_1044 VGND VPWR sky130_fd_sc_hd__fill_1
X_4564_ _4561_/X _4562_/X _4581_/A _4566_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_116_533 VGND VPWR sky130_fd_sc_hd__decap_12
X_6303_ _5978_/X _6073_/X _6302_/X _7750_/Q _6084_/X _6304_/B VGND VPWR sky130_fd_sc_hd__a32oi_4
X_7283_ _7282_/Y _7300_/B _7283_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4495_ _4495_/A _4495_/B _4495_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_116_566 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_886 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_428 VGND VPWR sky130_fd_sc_hd__decap_12
X_6234_ _6219_/A _6232_/X _6233_/X _5062_/A _6109_/X _6234_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_116_599 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1140 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_1102 VGND VPWR sky130_fd_sc_hd__decap_12
X_6165_ _5042_/X _6165_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_98_973 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1143 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1146 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_303 VGND VPWR sky130_fd_sc_hd__fill_2
X_5116_ _5107_/X _5113_/X _5114_/X _5115_/X _5116_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_100_934 VGND VPWR sky130_fd_sc_hd__decap_12
X_6096_ _6025_/X _4448_/X _6096_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_85_645 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_1187 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_196 VGND VPWR sky130_fd_sc_hd__decap_12
X_5047_ _5046_/X _5047_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_72_306 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_166 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_150_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_328 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_520 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_391 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6998_ _6932_/A la_data_in[76] _6934_/X _6998_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XPHY_3949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_266 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_558 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_428 VGND VPWR sky130_fd_sc_hd__decap_12
X_5949_ _5944_/X _5946_/Y _5947_/X _5948_/X _5949_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_209_1080 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_236 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_912 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1248 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_995 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1199 VGND VPWR sky130_fd_sc_hd__decap_3
X_7619_ _7139_/X _7619_/Q _7624_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_194_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_959 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_330 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1024 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_661 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_577 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_536 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_1079 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_794 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_1219 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_369 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_1151 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_520 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1093 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_350 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1077 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1107 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_288 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_250 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_900 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_261 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_962 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_731 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_283 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_294 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_977 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1050 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_704 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_1241 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_812 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_300 VGND VPWR sky130_fd_sc_hd__decap_12
X_4280_ _4276_/X _4279_/B _4279_/X _4280_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_180_491 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_818 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_881 VGND VPWR sky130_fd_sc_hd__decap_4
X_6921_ _6863_/X _6919_/X _6920_/Y _6921_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_81_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_851 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_542 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1212 VGND VPWR sky130_fd_sc_hd__decap_8
X_6852_ _7653_/Q _6852_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_63_873 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1245 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_895 VGND VPWR sky130_fd_sc_hd__decap_12
X_5803_ _5783_/X _5802_/X _5803_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_62_383 VGND VPWR sky130_fd_sc_hd__decap_12
X_6783_ _6767_/X _6781_/X _6782_/Y _6783_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_3995_ _3995_/A _6028_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_167_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_838 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_337 VGND VPWR sky130_fd_sc_hd__decap_8
X_5734_ _5731_/X _5732_/X _5733_/X _5734_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_206_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1128 VGND VPWR sky130_fd_sc_hd__fill_1
X_5665_ _5660_/X _5661_/X _5660_/X _5661_/X _5665_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_129_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_403 VGND VPWR sky130_fd_sc_hd__decap_12
X_7404_ _7404_/A _7404_/B _7403_/Y _7404_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_4616_ _4615_/A _4615_/B _4615_/X _4616_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_148_499 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_639 VGND VPWR sky130_fd_sc_hd__fill_2
X_5596_ _5594_/X _5595_/X _5593_/X _5597_/B VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_159_1038 VGND VPWR sky130_fd_sc_hd__decap_12
X_7335_ _7335_/A _7351_/B _7335_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_128_190 VGND VPWR sky130_fd_sc_hd__decap_12
X_4547_ _4547_/A _4590_/B _4549_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_132_801 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_992 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1257 VGND VPWR sky130_fd_sc_hd__decap_12
X_7266_ _7263_/Y _7265_/X _7266_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_143_171 VGND VPWR sky130_fd_sc_hd__decap_12
X_4478_ _4820_/B _4479_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_116_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_867 VGND VPWR sky130_fd_sc_hd__fill_1
X_6217_ _4794_/Y _6216_/X _6194_/X _6217_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_89_269 VGND VPWR sky130_fd_sc_hd__decap_12
X_7197_ _7224_/A _7224_/B _7225_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_86_910 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_921 VGND VPWR sky130_fd_sc_hd__decap_12
X_6148_ _6148_/A _6011_/X _6149_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_161_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_591 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_678 VGND VPWR sky130_fd_sc_hd__decap_12
X_6079_ _6027_/Y _6028_/B _4036_/A _6079_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_161_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_1028 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_177 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_22_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_300 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_873 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_715 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_4469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_501 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_681 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_79 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_534 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_849 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_580 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_229 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_753 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_925 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_820 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_864 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_970 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_672 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_108_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_867 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_718 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_910 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1032 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_623 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1212 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_114_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_818 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_328 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_445 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_810 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_394 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_517 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_556 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_90 VGND VPWR sky130_fd_sc_hd__fill_2
X_3780_ _4769_/A _4552_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_73_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_898 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1142 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_509 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_550 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_893 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_263 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_785 VGND VPWR sky130_fd_sc_hd__decap_8
X_5450_ _5446_/Y _5449_/X _5446_/Y _5449_/X _5450_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_157_285 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_959 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_756 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_4401_ _4400_/A _4400_/B _4400_/X _4401_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_201_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_650 VGND VPWR sky130_fd_sc_hd__decap_3
X_5381_ _5368_/X _5371_/X _5381_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_7120_ _7128_/A _7120_/B _7120_/C _7626_/D VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_160_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_288 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_2_0_wb_clk_i clkbuf_3_3_0_wb_clk_i/A clkbuf_3_2_0_wb_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4332_ _4331_/A _4331_/B _4331_/X _4332_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_119_1011 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_62 VGND VPWR sky130_fd_sc_hd__decap_12
X_7051_ _7049_/Y _7050_/Y _7049_/Y _7050_/Y _7117_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_141_664 VGND VPWR sky130_fd_sc_hd__decap_6
X_4263_ _4554_/A _4394_/B _4263_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_140_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_517 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1088 VGND VPWR sky130_fd_sc_hd__decap_8
X_6002_ _5573_/Y _5574_/Y _6002_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_119_1099 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_239 VGND VPWR sky130_fd_sc_hd__decap_12
X_4194_ _4156_/X _4193_/X _4156_/X _4193_/X _4194_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_83_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_464 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_998 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_626 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_434 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1001 VGND VPWR sky130_fd_sc_hd__decap_12
X_6904_ _6840_/A la_data_in[55] _6842_/X _6904_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_70_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_501 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_602 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1004 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_1056 VGND VPWR sky130_fd_sc_hd__fill_1
X_6835_ la_data_in[57] _6835_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_196_815 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_1078 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_837 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1048 VGND VPWR sky130_fd_sc_hd__decap_8
X_6766_ _6723_/A _6723_/B _6723_/X _6765_/X _6766_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XPHY_1629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1059 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_729 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_206 VGND VPWR sky130_fd_sc_hd__decap_8
X_3978_ _3976_/X _3977_/X _3975_/X _3978_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_52_1223 VGND VPWR sky130_fd_sc_hd__decap_8
X_5717_ _5704_/X _5705_/X _5715_/X _5716_/X _5717_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_210_178 VGND VPWR sky130_fd_sc_hd__decap_12
X_6697_ _6647_/A _6647_/B _6697_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_109_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_15 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_5648_ _5492_/X _5493_/X _5492_/X _5493_/X _5648_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_164_745 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_447 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_469 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_650 VGND VPWR sky130_fd_sc_hd__decap_12
X_5579_ _5579_/A _5578_/X _5580_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_117_672 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_1081 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_428 VGND VPWR sky130_fd_sc_hd__decap_12
X_7318_ _4747_/A _7293_/X _7317_/X _7318_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_105_834 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1005 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_355 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_1038 VGND VPWR sky130_fd_sc_hd__decap_12
X_7249_ wbs_cyc_i wbs_stb_i _7238_/A _7249_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_120_837 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_818 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_998 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_572 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_1121 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_171_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_147 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1093 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1112 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1240 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_670 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_361 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_117 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_62 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1153 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1156 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_4299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1186 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_567 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_123 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_364 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_70 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1252 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_962 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_950 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1146 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_526 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_848 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_994 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_212 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_467 VGND VPWR sky130_fd_sc_hd__decap_3
X_4950_ _7773_/Q _4900_/B _5023_/B _4950_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_80_938 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_440 VGND VPWR sky130_fd_sc_hd__decap_12
X_3901_ _3900_/Y _3901_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_75_1245 VGND VPWR sky130_fd_sc_hd__decap_6
X_4881_ _4881_/A _4881_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_178_837 VGND VPWR sky130_fd_sc_hd__decap_12
X_6620_ _6618_/Y _6619_/Y _6618_/Y _6619_/Y _6620_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_3832_ _3832_/A _3832_/B _3832_/C _3832_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_189_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_818 VGND VPWR sky130_fd_sc_hd__decap_12
X_6551_ _6500_/A _6500_/B _6500_/X _6550_/X _6551_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_3763_ _3763_/A _4570_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_203_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_572 VGND VPWR sky130_fd_sc_hd__decap_8
X_5502_ _4467_/A _5275_/X _5502_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_199_1160 VGND VPWR sky130_fd_sc_hd__decap_12
X_6482_ _6427_/X _6479_/X _6481_/X _6482_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_3694_ wbs_adr_i[1] wbs_adr_i[0] wbs_adr_i[3] wbs_adr_i[2] _3710_/A VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_195_1013 VGND VPWR sky130_fd_sc_hd__decap_12
X_5433_ _5419_/X _5425_/X _5419_/X _5425_/X _5433_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_69_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1046 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_417 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_156_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_428 VGND VPWR sky130_fd_sc_hd__decap_12
X_5364_ _5363_/A _5363_/B _5363_/X _5364_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_99_342 VGND VPWR sky130_fd_sc_hd__decap_12
X_7103_ _7128_/A _7095_/X _7102_/Y _7103_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_4315_ _4255_/X _4313_/X _4310_/X _4314_/X _4315_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_102_815 VGND VPWR sky130_fd_sc_hd__decap_8
X_5295_ _5293_/X _5294_/X _5293_/X _5294_/X _5295_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_59_228 VGND VPWR sky130_fd_sc_hd__decap_12
X_7034_ _7034_/A _7034_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4246_ _4240_/X _4241_/X _4239_/X _4242_/X _4246_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_102_859 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_902 VGND VPWR sky130_fd_sc_hd__decap_8
X_4177_ _4157_/X _4176_/X _4157_/X _4176_/X _4177_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_210_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1052 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_870 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_570 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_607 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_15 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_489 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_459 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1167 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_364 VGND VPWR sky130_fd_sc_hd__fill_2
X_6818_ _6912_/A _6814_/A _6817_/X _7666_/D VGND VPWR sky130_fd_sc_hd__and3_4
XPHY_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_898 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7798_ _7798_/D _3867_/A _7801_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_1020 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1140 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_537 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_550 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1042 VGND VPWR sky130_fd_sc_hd__decap_12
X_6749_ la_data_in[33] _6749_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_17_1184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_288 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_279 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_1160 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1250 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_1182 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_710 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1166 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_207_716 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_423 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1185 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_776 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_32 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_640 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_410 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_70 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_971 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_81 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_92 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_673 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1243 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_840 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1137 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_756 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_80 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_361 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_970 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_726 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_992 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_556 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_247 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_1022 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_802 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_995 VGND VPWR sky130_fd_sc_hd__decap_12
X_4100_ _4098_/X _4099_/X _4101_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_151_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_334 VGND VPWR sky130_fd_sc_hd__fill_2
X_5080_ _4666_/A _4915_/B _5080_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_155_1096 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_645 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_41 VGND VPWR sky130_fd_sc_hd__decap_8
X_4031_ _4026_/X _4028_/X _4029_/Y _4030_/X _4031_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_110_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_52 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_401 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_434 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_456 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_916 VGND VPWR sky130_fd_sc_hd__decap_12
X_5982_ _5941_/X _5942_/X _5941_/X _5942_/X _6293_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_37_489 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_52_437 VGND VPWR sky130_fd_sc_hd__decap_12
X_4933_ _4865_/X _4866_/X _4859_/X _4867_/X _4933_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_7721_ _6471_/X _7721_/Q _7785_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_205_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1015 VGND VPWR sky130_fd_sc_hd__decap_12
X_4864_ _4861_/X _4863_/B _4863_/X _4864_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_7652_ _6921_/X _7652_/Q _7758_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_33_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1097 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_807 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_13 _6190_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_178_678 VGND VPWR sky130_fd_sc_hd__decap_12
X_3815_ wbs_dat_i[11] _3822_/B _3815_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_6603_ _7695_/Q _6605_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_7583_ _7583_/HI la_data_out[110] VGND VPWR sky130_fd_sc_hd__conb_1
X_4795_ _4792_/X _4793_/X _4792_/X _4793_/X _4795_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6534_ _6531_/Y _6532_/Y _6531_/Y _6532_/Y _6596_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_520 VGND VPWR sky130_fd_sc_hd__decap_8
X_3746_ _4485_/A _4919_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_193_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_745 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_767 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1086 VGND VPWR sky130_fd_sc_hd__decap_12
X_6465_ _6057_/A _6465_/B _6464_/Y _7723_/D VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_161_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_5416_ _5407_/X _5415_/X _5407_/X _5415_/X _5416_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_173_394 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_940 VGND VPWR sky130_fd_sc_hd__decap_4
X_6396_ _6396_/A _6396_/B _6396_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_88_802 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1182 VGND VPWR sky130_fd_sc_hd__decap_8
X_5347_ _5137_/A _4756_/B _5347_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_114_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_943 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_857 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_954 VGND VPWR sky130_fd_sc_hd__decap_12
X_5278_ _5274_/X _5276_/X _5274_/X _5276_/X _5278_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_102_667 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_367 VGND VPWR sky130_fd_sc_hd__decap_12
X_7017_ _6976_/X _7016_/X _6999_/X _7017_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_4229_ _3738_/A _4546_/B _4229_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_28_412 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_1024 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_581 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_404 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_724 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_938 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_601 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_971 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_150 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1159 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_818 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_273 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_200_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_317 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_367 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1041 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_810 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_726 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_832 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1036 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_556 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_802 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_566 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_1203 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_835 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_483 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_312 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_431 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_987 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_849 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_497 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1031 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1192 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_489 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_1034 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_212 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1059 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_448 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_420 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_3170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_684 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_453 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_785 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_306 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_520 VGND VPWR sky130_fd_sc_hd__decap_12
X_4580_ _4580_/A _4580_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_1790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_862 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_1130 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_821 VGND VPWR sky130_fd_sc_hd__decap_12
X_6250_ _5778_/X _6249_/X _6250_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_66_1008 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_331 VGND VPWR sky130_fd_sc_hd__decap_4
X_5201_ _5199_/X _5201_/B _5201_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_157_1158 VGND VPWR sky130_fd_sc_hd__fill_1
X_6181_ _4949_/A _6158_/X _6144_/X _6181_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_124_770 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_910 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_386 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_921 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_239 VGND VPWR sky130_fd_sc_hd__decap_12
X_5132_ _5129_/X _5130_/X _5131_/X _5132_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_69_367 VGND VPWR sky130_fd_sc_hd__decap_12
X_5063_ _4513_/A _4479_/B _5063_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_84_337 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1052 VGND VPWR sky130_fd_sc_hd__decap_12
X_4014_ _4535_/A _4123_/B _4014_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_37_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_562 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_297 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_1276 VGND VPWR sky130_fd_sc_hd__fill_1
X_5965_ _5200_/A _4491_/A _5972_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_52_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_407 VGND VPWR sky130_fd_sc_hd__decap_12
X_7704_ _6584_/X _7704_/Q _7696_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4916_ _4570_/A _4844_/B _4916_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_5896_ _5892_/X _5893_/X _5894_/Y _5895_/X _5896_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_139_818 VGND VPWR sky130_fd_sc_hd__decap_12
X_7635_ _7031_/X _6965_/A _7624_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_178_475 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_4847_ _4847_/A _4847_/B _4847_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_138_317 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_637 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_4778_ _4498_/A _4778_/B _4779_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7566_ _7566_/HI la_data_out[93] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_165_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_478 VGND VPWR sky130_fd_sc_hd__decap_8
X_3729_ _3728_/X _4494_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_6517_ la_data_in[6] _6518_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_193_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_884 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_146_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_895 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_586 VGND VPWR sky130_fd_sc_hd__decap_12
X_7497_ _7497_/HI la_data_out[24] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_162_832 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1217 VGND VPWR sky130_fd_sc_hd__decap_3
X_6448_ _6381_/A _6446_/Y _6448_/C _6448_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_164_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_718 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_898 VGND VPWR sky130_fd_sc_hd__fill_2
X_6379_ _5275_/X _6345_/A _6381_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_0_525 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_965 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_453 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_816 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_507 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_529 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1130 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_795 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_348 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1174 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_242 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1204 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1219 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1218 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_245 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_459 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_410 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_421 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_289 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_632 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1062 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_306 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_974 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_755 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_996 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_659 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_788 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_146 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_873 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_523 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_820 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_843 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1063 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1044 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1006 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1069 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1129 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_170_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_286 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_234 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_418 VGND VPWR sky130_fd_sc_hd__decap_3
X_5750_ _4747_/A _5533_/B _5750_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_50_738 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_740 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1102 VGND VPWR sky130_fd_sc_hd__fill_1
X_4701_ _4546_/X _4550_/X _4546_/X _4550_/X _4701_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_5681_ _5348_/A _4363_/A _5681_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_198_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1089 VGND VPWR sky130_fd_sc_hd__fill_2
X_4632_ _3771_/A _4277_/A _4634_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_7420_ io_oeb[15] _7420_/LO VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_147_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_873 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_84 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_489 VGND VPWR sky130_fd_sc_hd__decap_12
X_4563_ _4561_/X _4562_/X _4581_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_7351_ _7351_/A _7351_/B _7351_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_162_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_990 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_426 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_821 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_1067 VGND VPWR sky130_fd_sc_hd__fill_1
X_6302_ _6299_/Y _6300_/Y _6301_/Y _6302_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_143_320 VGND VPWR sky130_fd_sc_hd__decap_12
X_7282_ io_in[9] _7282_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_190_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_545 VGND VPWR sky130_fd_sc_hd__fill_2
X_4494_ _4494_/A _4493_/X _4495_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_6_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_407 VGND VPWR sky130_fd_sc_hd__decap_12
X_6233_ _6223_/Y _6225_/Y _6233_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_116_589 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_397 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1152 VGND VPWR sky130_fd_sc_hd__decap_6
X_6164_ _6185_/A _6164_/B _7776_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_44_1114 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_985 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_462 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_1196 VGND VPWR sky130_fd_sc_hd__decap_12
X_5115_ _5107_/X _5113_/X _5107_/X _5113_/X _5115_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_170_1155 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1158 VGND VPWR sky130_fd_sc_hd__decap_8
X_6095_ _6095_/A _6095_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_5046_ _5045_/X _5046_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_211_1141 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_679 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_178 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_532 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_504 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1013 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1241 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6997_ _6985_/X _6995_/X _6996_/Y _6997_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_20_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1057 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_278 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1221 VGND VPWR sky130_fd_sc_hd__decap_12
X_5948_ _5913_/X _5917_/X _5913_/X _5917_/X _5948_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_159_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_941 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_1092 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_248 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_615 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_440 VGND VPWR sky130_fd_sc_hd__decap_12
X_5879_ _5850_/X _5851_/X _5850_/X _5851_/X _5879_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_159_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_473 VGND VPWR sky130_fd_sc_hd__decap_12
X_7618_ _7141_/X _7618_/Q _7624_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_194_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_501 VGND VPWR sky130_fd_sc_hd__decap_8
X_7549_ _7549_/HI la_data_out[76] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_135_821 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_1090 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_448 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_1036 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_971 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_673 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_801 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_175_1055 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_589 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_812 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_823 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_846 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1203 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_619 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_871 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_562 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1061 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_1196 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_1038 VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_4_0_wb_clk_i clkbuf_3_2_0_wb_clk_i/X _7696_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_17_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1004 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_204_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_82 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_147_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1026 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1089 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_1119 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_749 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_240 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_251 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_912 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_273 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_974 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_284 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_295 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_489 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_865 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_661 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_684 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1237 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_315 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_977 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_178 VGND VPWR sky130_fd_sc_hd__decap_12
X_6920_ _6863_/X _6919_/X _6905_/X _6920_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_81_159 VGND VPWR sky130_fd_sc_hd__decap_12
X_6851_ _6849_/Y _6850_/Y _6849_/Y _6850_/Y _6866_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_207_184 VGND VPWR sky130_fd_sc_hd__decap_12
X_5802_ _5784_/X _5801_/B _5801_/X _5802_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_22_215 VGND VPWR sky130_fd_sc_hd__decap_4
X_3994_ _3994_/A _3993_/Y _3995_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_6782_ _6767_/X _6781_/X _6690_/X _6782_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_62_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_149_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_557 VGND VPWR sky130_fd_sc_hd__fill_1
X_5733_ _5731_/X _5732_/X _5733_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_188_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_771 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_220 VGND VPWR sky130_fd_sc_hd__decap_12
X_5664_ _5654_/X _5663_/X _5654_/X _5663_/X _5664_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_176_776 VGND VPWR sky130_fd_sc_hd__decap_12
X_7403_ wbs_dat_i[24] _3882_/X _7403_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_4615_ _4615_/A _4615_/B _4615_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_163_415 VGND VPWR sky130_fd_sc_hd__decap_12
X_5595_ _5198_/A _4631_/B _5595_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_159_1028 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_40 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_62 VGND VPWR sky130_fd_sc_hd__decap_8
X_4546_ _4645_/A _4546_/B _4546_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7334_ _7276_/A _7351_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_102_1274 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_813 VGND VPWR sky130_fd_sc_hd__decap_8
X_4477_ _4477_/A _4820_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_7265_ _7276_/A _7265_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_145_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1269 VGND VPWR sky130_fd_sc_hd__decap_8
X_6216_ _6317_/C _6216_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_7196_ _7160_/Y _7161_/Y _7227_/B _7224_/B VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_135_1050 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_6147_ _5032_/B _6147_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_112_581 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_944 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_161_27 VGND VPWR sky130_fd_sc_hd__decap_12
X_6078_ _6028_/A _6081_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_100_776 VGND VPWR sky130_fd_sc_hd__fill_2
X_5029_ _5017_/X _5026_/X _5027_/X _5028_/X _5029_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XPHY_4404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_690 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_351 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_69 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_693 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_568 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_900 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1032 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_1095 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_765 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_944 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_1016 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_618 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1038 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_937 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_999 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_832 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_876 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_813 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_108_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_790 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_846 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_345 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_602 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_675 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1236 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_686 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_646 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1258 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_903 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_167 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_947 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_457 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_576 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_529 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1168 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_584 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_297 VGND VPWR sky130_fd_sc_hd__decap_8
X_4400_ _4400_/A _4400_/B _4400_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_173_768 VGND VPWR sky130_fd_sc_hd__fill_1
X_5380_ _5337_/X _5358_/X _5378_/X _5379_/X _5380_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_201_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_971 VGND VPWR sky130_fd_sc_hd__decap_12
X_4331_ _4331_/A _4331_/B _4331_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_5_74 VGND VPWR sky130_fd_sc_hd__decap_12
X_7050_ la_data_in[89] _7050_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4262_ _4514_/A _4217_/B _4264_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_99_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_367 VGND VPWR sky130_fd_sc_hd__decap_12
X_6001_ _5548_/X _5564_/X _6011_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_101_529 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_922 VGND VPWR sky130_fd_sc_hd__fill_1
X_4193_ _4157_/X _4176_/X _4177_/X _4192_/X _4193_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_68_944 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_471 VGND VPWR sky130_fd_sc_hd__decap_12
X_6903_ _6912_/A _6872_/X _6903_/C _6903_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_165_1010 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_660 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_1013 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_513 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_63 VGND VPWR sky130_fd_sc_hd__decap_12
X_6834_ _6834_/A _6834_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_211_614 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_321 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_855 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_168_518 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_849 VGND VPWR sky130_fd_sc_hd__decap_6
X_6765_ _6724_/Y _6725_/Y _6764_/X _6765_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_91_1262 VGND VPWR sky130_fd_sc_hd__decap_12
X_3977_ _3722_/A _4164_/B _3977_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_50_376 VGND VPWR sky130_fd_sc_hd__decap_12
X_5716_ _5704_/X _5705_/X _5704_/X _5705_/X _5716_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_176_540 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_1208 VGND VPWR sky130_fd_sc_hd__decap_12
X_6696_ _6694_/X _6696_/B _6696_/C _6696_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_137_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_629 VGND VPWR sky130_fd_sc_hd__decap_12
X_5647_ _5645_/X _5646_/X _5647_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_108_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_459 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_919 VGND VPWR sky130_fd_sc_hd__decap_8
X_5578_ _5328_/X _5329_/X _5289_/X _5330_/X _5578_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_117_662 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_587 VGND VPWR sky130_fd_sc_hd__decap_12
X_7317_ _7316_/Y _7324_/B _7317_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_176_1150 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_684 VGND VPWR sky130_fd_sc_hd__decap_12
X_4529_ _7769_/Q _4529_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_105_846 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_323 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_952 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_654 VGND VPWR sky130_fd_sc_hd__decap_12
X_7248_ _7238_/A _7245_/A _7247_/X _7602_/D VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_105_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_410 VGND VPWR sky130_fd_sc_hd__decap_12
X_7179_ la_data_in[98] _7180_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_46_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_413 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_947 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_159 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_811 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1124 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_682 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_129 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_74 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_192 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1059 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_579 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_135 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_220 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_590 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_871 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_712 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_919 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_727 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_470 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_82 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_1275 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_708 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_985 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_1158 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_473 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_687 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_202 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_224 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_115 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1161 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_852 VGND VPWR sky130_fd_sc_hd__decap_12
X_3900_ _6319_/A _3900_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_205_452 VGND VPWR sky130_fd_sc_hd__decap_12
X_4880_ _4809_/X _4879_/X _4809_/X _4879_/X _4880_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_33_855 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1227 VGND VPWR sky130_fd_sc_hd__decap_12
X_3831_ wbs_dat_i[9] _3822_/B _3832_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_178_849 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_398 VGND VPWR sky130_fd_sc_hd__decap_12
X_3762_ _7811_/Q _3763_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_6550_ _6503_/A _6502_/Y _6503_/X _6549_/X _6550_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_119_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1082 VGND VPWR sky130_fd_sc_hd__fill_1
X_5501_ _5501_/A _5491_/X _5501_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_203_1257 VGND VPWR sky130_fd_sc_hd__decap_12
X_3693_ _4535_/A _3693_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_6481_ _6670_/A _6481_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_185_381 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_459 VGND VPWR sky130_fd_sc_hd__decap_12
X_5432_ _5431_/A _5430_/X _5431_/X _5432_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_195_1025 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_779 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1252 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_5363_ _5363_/A _5363_/B _5363_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_154_790 VGND VPWR sky130_fd_sc_hd__decap_8
X_7102_ _7095_/A _7095_/B _7102_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_4314_ _4255_/X _4313_/X _4255_/X _4313_/X _4314_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_354 VGND VPWR sky130_fd_sc_hd__decap_12
X_5294_ _5294_/A _5294_/B _5294_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_99_387 VGND VPWR sky130_fd_sc_hd__fill_2
X_4245_ _4214_/X _4244_/X _4214_/X _4244_/X _4245_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7033_ _7012_/A _7030_/A _7032_/X _7634_/D VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_45_1050 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_741 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_4176_ _4158_/X _4165_/X _4166_/X _4175_/X _4176_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_132_1064 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_882 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_733 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1138 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_619 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_276 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_304 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6817_ _7666_/Q la_data_in[32] _6817_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_2139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7797_ _7797_/D _3875_/A _7797_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_337 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1179 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_359 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_466 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_398 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1100 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1081 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_1152 VGND VPWR sky130_fd_sc_hd__decap_6
X_6748_ _6748_/A _6748_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_167_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_871 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1054 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_724 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_595 VGND VPWR sky130_fd_sc_hd__decap_12
X_6679_ _6612_/A la_data_in[26] _6614_/X _6679_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_164_532 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_746 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_971 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_727 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_481 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_613 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_240 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_1142 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_1194 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_785 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_882 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_722 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_958 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_728 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_295 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_435 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1189 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_227 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_405 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_811 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_44 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_912 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_440 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_855 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_60 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_202_422 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_82 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_983 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_93 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_685 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_825 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1110 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_184 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_858 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1154 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1187 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_1149 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_571 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_852 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_407 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_941 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1061 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1034 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_1106 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_814 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_602 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_1037 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_657 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1212 VGND VPWR sky130_fd_sc_hd__decap_12
X_4030_ _4026_/X _4028_/X _4026_/X _4028_/X _4030_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_64 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_413 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_733 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_468 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_714 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_928 VGND VPWR sky130_fd_sc_hd__decap_12
X_5981_ _5950_/X _5952_/X _5980_/X _5983_/A VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_64_276 VGND VPWR sky130_fd_sc_hd__decap_12
X_7720_ _6474_/X _7720_/Q _7785_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4932_ _4928_/X _4931_/X _4928_/X _4931_/X _4932_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_52_449 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_1111 VGND VPWR sky130_fd_sc_hd__decap_12
X_7651_ _7651_/D _7651_/Q _7756_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_205_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1027 VGND VPWR sky130_fd_sc_hd__decap_4
X_4863_ _4861_/X _4863_/B _4863_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_177_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_471 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_696 VGND VPWR sky130_fd_sc_hd__decap_12
X_6602_ _6600_/Y _6601_/Y _6600_/Y _6601_/Y _6602_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_123_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_14 _7263_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_3814_ _3813_/X _3798_/B _3814_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_166_819 VGND VPWR sky130_fd_sc_hd__decap_4
X_7582_ _7582_/HI la_data_out[109] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_335 VGND VPWR sky130_fd_sc_hd__fill_1
X_4794_ _7767_/Q _4794_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_6533_ _7698_/Q la_data_in[0] _6596_/A VGND VPWR sky130_fd_sc_hd__nand2_4
X_3745_ _4613_/A _4485_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_186_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_779 VGND VPWR sky130_fd_sc_hd__decap_12
X_6464_ _6399_/X _6464_/B _6464_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_134_716 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_727 VGND VPWR sky130_fd_sc_hd__decap_12
X_5415_ _5413_/X _5414_/X _5413_/X _5414_/X _5415_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6395_ la_data_in[122] _6396_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_12_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1123 VGND VPWR sky130_fd_sc_hd__decap_12
X_5346_ _5339_/X _5345_/X _5346_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_88_814 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_911 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1009 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_495 VGND VPWR sky130_fd_sc_hd__decap_12
X_5277_ _7762_/Q _5277_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_101_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_966 VGND VPWR sky130_fd_sc_hd__decap_12
X_7016_ _6950_/A la_data_in[70] _6952_/X _7016_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_4228_ _4624_/B _4546_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_87_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_4159_ _4499_/A _4217_/B _4162_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_210_1036 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_619 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_107 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1252 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1271 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_1105 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_983 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_162 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_825 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_836 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_184 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_605 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_306 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_329 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1020 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_874 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1053 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_844 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_847 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_944 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_966 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_443 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_977 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_999 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_891 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1160 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1043 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_928 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_1076 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1008 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_224 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_257 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_944 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_199_281 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_696 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_263 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_318 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_80 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_80 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_833 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_855 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_866 VGND VPWR sky130_fd_sc_hd__decap_12
X_5200_ _5200_/A _4648_/A _5201_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_131_719 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3 VGND VPWR sky130_fd_sc_hd__decap_8
X_6180_ _4983_/X _6178_/X _6101_/X _6180_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_97_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_933 VGND VPWR sky130_fd_sc_hd__decap_12
X_5131_ _5129_/X _5130_/X _5131_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_123_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_806 VGND VPWR sky130_fd_sc_hd__decap_12
X_5062_ _5062_/A _5062_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_96_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_379 VGND VPWR sky130_fd_sc_hd__decap_6
X_4013_ _4006_/X _4012_/X _4006_/X _4012_/X _4013_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_722 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1064 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1211 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_86 VGND VPWR sky130_fd_sc_hd__decap_12
X_5964_ _5959_/X _5960_/X _5959_/X _5960_/X _5974_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_52_257 VGND VPWR sky130_fd_sc_hd__fill_1
X_7703_ _6586_/X _7703_/Q _7696_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_178_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_577 VGND VPWR sky130_fd_sc_hd__decap_3
X_4915_ _4519_/A _4915_/B _4915_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_40_419 VGND VPWR sky130_fd_sc_hd__decap_12
X_5895_ _5892_/X _5893_/X _5892_/X _5893_/X _5895_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_21_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_977 VGND VPWR sky130_fd_sc_hd__decap_8
X_7634_ _7634_/D _6967_/A _7624_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_178_465 VGND VPWR sky130_fd_sc_hd__fill_1
X_4846_ _4842_/X _4844_/X _4845_/X _4846_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_178_487 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_329 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_53_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_649 VGND VPWR sky130_fd_sc_hd__decap_12
X_7565_ _7565_/HI la_data_out[92] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_140_1130 VGND VPWR sky130_fd_sc_hd__decap_12
X_4777_ _4562_/B _4778_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_165_159 VGND VPWR sky130_fd_sc_hd__decap_12
X_6516_ _7704_/Q _6516_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_14_1166 VGND VPWR sky130_fd_sc_hd__decap_12
X_3728_ _4561_/A _3728_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_10_1008 VGND VPWR sky130_fd_sc_hd__decap_12
X_7496_ _7496_/HI la_data_out[23] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_174_671 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1158 VGND VPWR sky130_fd_sc_hd__fill_1
X_6447_ la_data_in[127] _6447_/B _6448_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_162_844 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_134_579 VGND VPWR sky130_fd_sc_hd__fill_1
X_6378_ _6381_/A _6378_/B _6377_/Y _7731_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_115_771 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_110 VGND VPWR sky130_fd_sc_hd__decap_12
X_5329_ _5211_/X _5226_/X _5120_/X _5227_/X _5329_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_138_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_559 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_839 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1115 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_541 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1186 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_703 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_777 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1216 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_883 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_86 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_400 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1060 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_411 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_410 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_422 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_471 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_903 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_110 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_465 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1074 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_318 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_424 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_457 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_158 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_395 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_535 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_708 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_579 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1170 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_741 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_1075 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_806 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_785 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1018 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_349 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_208_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_845 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_769 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_246 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_550 VGND VPWR sky130_fd_sc_hd__decap_4
X_4700_ _4695_/X _4699_/X _4698_/X _4700_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_176_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_605 VGND VPWR sky130_fd_sc_hd__decap_12
X_5680_ _5615_/X _5619_/X _5615_/X _5619_/X _5680_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_72_1057 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_964 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_947 VGND VPWR sky130_fd_sc_hd__decap_8
X_4631_ _4503_/A _4631_/B _4631_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_198_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_969 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_147_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_863 VGND VPWR sky130_fd_sc_hd__decap_3
X_7350_ io_in[21] _7351_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_163_619 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_928 VGND VPWR sky130_fd_sc_hd__decap_12
X_4562_ _4479_/A _4562_/B _4562_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_129_885 VGND VPWR sky130_fd_sc_hd__decap_4
X_6301_ _5954_/X _5963_/X _5954_/X _5963_/X _6301_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_156_693 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_7281_ _7781_/Q _7260_/B _7281_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_7_692 VGND VPWR sky130_fd_sc_hd__fill_1
X_4493_ _4565_/B _4493_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_6232_ _6223_/A _6225_/A _6232_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_89_419 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1101 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_110 VGND VPWR sky130_fd_sc_hd__decap_12
X_6163_ _6106_/X _6161_/X _6162_/X _4434_/A _6109_/X _6164_/B VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_44_1126 VGND VPWR sky130_fd_sc_hd__decap_3
X_5114_ _5055_/X _5056_/X _5055_/X _5056_/X _5114_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_85_603 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_997 VGND VPWR sky130_fd_sc_hd__decap_8
X_6094_ _6089_/X _6090_/X _6093_/X _6094_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_170_1167 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_796 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_284 VGND VPWR sky130_fd_sc_hd__decap_12
X_5045_ _5045_/A _5045_/B _5045_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_66_861 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_842 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_516 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_1025 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1170 VGND VPWR sky130_fd_sc_hd__fill_1
X_6996_ _6985_/X _6995_/X _6905_/X _6996_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XPHY_3929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1253 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1200 VGND VPWR sky130_fd_sc_hd__decap_12
X_5947_ _5944_/X _5946_/Y _5944_/X _5946_/Y _5947_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_129_1069 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_251 VGND VPWR sky130_fd_sc_hd__decap_12
X_5878_ _5859_/X _5878_/B _5878_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_179_785 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_452 VGND VPWR sky130_fd_sc_hd__decap_6
X_7617_ _7617_/D io_out[6] _7797_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4829_ _4829_/A _4613_/B _4829_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_193_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_485 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_166_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_788 VGND VPWR sky130_fd_sc_hd__decap_12
X_7548_ _7548_/HI la_data_out[75] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_175_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_844 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_630 VGND VPWR sky130_fd_sc_hd__decap_8
X_7479_ _7479_/HI la_data_out[6] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_175_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_855 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_983 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_931 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_356 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_541 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_883 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_382 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_596 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_50 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_886 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_147_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_230 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_252 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_750 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_520 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_274 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_733 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_60 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_285 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_71 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_811 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_877 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_1265 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1145 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_673 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1249 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_485 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_327 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_308 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_664 VGND VPWR sky130_fd_sc_hd__decap_12
X_6850_ la_data_in[52] _6850_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_74_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_566 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_196 VGND VPWR sky130_fd_sc_hd__decap_12
X_5801_ _5784_/X _5801_/B _5801_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_211_807 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_205 VGND VPWR sky130_fd_sc_hd__decap_8
X_6781_ _6715_/A la_data_in[44] _6717_/X _6781_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_3993_ _3993_/A _3991_/X _3993_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_200_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_317 VGND VPWR sky130_fd_sc_hd__decap_12
X_5732_ _5186_/A _4291_/A _5732_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_176_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_249 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_958 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_783 VGND VPWR sky130_fd_sc_hd__decap_8
X_5663_ _5655_/X _5662_/X _5655_/X _5662_/X _5663_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_148_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1130 VGND VPWR sky130_fd_sc_hd__decap_8
X_7402_ _3918_/X _3897_/B _7404_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_191_703 VGND VPWR sky130_fd_sc_hd__decap_12
X_4614_ _4614_/A _4830_/B _4615_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_176_788 VGND VPWR sky130_fd_sc_hd__decap_12
X_5594_ _5591_/X _5592_/X _5593_/X _5594_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_190_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1067 VGND VPWR sky130_fd_sc_hd__fill_1
X_7333_ io_in[18] _7335_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_209_52 VGND VPWR sky130_fd_sc_hd__decap_8
X_4545_ _4530_/X _4535_/X _4529_/Y _4536_/X _4545_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_117_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_74 VGND VPWR sky130_fd_sc_hd__decap_12
X_7264_ _7264_/A _7264_/B _7276_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_132_825 VGND VPWR sky130_fd_sc_hd__decap_12
X_4476_ _4475_/Y _4477_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_171_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_398 VGND VPWR sky130_fd_sc_hd__decap_8
X_6215_ _6212_/Y _6213_/X _6319_/C _6215_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_7195_ _7226_/A _7194_/X _7227_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_48_1081 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_379 VGND VPWR sky130_fd_sc_hd__decap_8
X_6146_ _6089_/X _6143_/X _6145_/X _6146_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_100_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_711 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_967 VGND VPWR sky130_fd_sc_hd__fill_1
X_6077_ _6308_/B _6189_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_161_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1008 VGND VPWR sky130_fd_sc_hd__fill_1
X_5028_ _5017_/X _5026_/X _5017_/X _5026_/X _5028_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_72_105 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_544 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_672 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_363 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6979_ _6946_/X _6978_/X _7012_/B VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_3759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1030 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_1000 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1052 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_1063 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_733 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_912 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_703 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_714 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_427 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_844 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_120 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_135_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_699 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_794 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_164 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1176 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_658 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_179 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_469 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_588 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_374 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1250 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_761 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_755 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_1196 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_777 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_503 VGND VPWR sky130_fd_sc_hd__decap_8
X_4330_ _4461_/A _4394_/B _4331_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_154_983 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_611 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1084 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1046 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_86 VGND VPWR sky130_fd_sc_hd__decap_12
X_4261_ _3786_/A _4514_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_45_1221 VGND VPWR sky130_fd_sc_hd__decap_12
X_6000_ _6008_/A _6000_/B _5584_/X _6000_/D _6148_/A VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_140_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_379 VGND VPWR sky130_fd_sc_hd__decap_12
X_4192_ _4186_/X _4191_/X _4186_/X _4191_/X _4192_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_95_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_444 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_135 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_1189 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_477 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_6902_ _6872_/A _6871_/X _6903_/C VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_35_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1180 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_970 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1022 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1025 VGND VPWR sky130_fd_sc_hd__decap_12
X_6833_ _6833_/A _6832_/Y _6833_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_78_1085 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_75 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1066 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_333 VGND VPWR sky130_fd_sc_hd__decap_3
X_6764_ _6792_/A _6763_/X _6764_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_1609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1039 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_709 VGND VPWR sky130_fd_sc_hd__decap_12
X_3976_ _3973_/X _3974_/X _3975_/X _3976_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_165_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1203 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1274 VGND VPWR sky130_fd_sc_hd__decap_3
X_5715_ _5711_/Y _5714_/X _5711_/Y _5714_/X _5715_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_50_388 VGND VPWR sky130_fd_sc_hd__decap_8
X_6695_ _6695_/A _6695_/B _6696_/C VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_164_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_928 VGND VPWR sky130_fd_sc_hd__decap_12
X_5646_ _5588_/X _5589_/X _5587_/X _5646_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_148_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_5577_ _5569_/X _5570_/X _5569_/X _5570_/X _5579_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_3_908 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_257 VGND VPWR sky130_fd_sc_hd__decap_12
X_7316_ io_in[15] _7316_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4528_ _4474_/X _4510_/X _4526_/X _4527_/X _4528_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_191_599 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_1094 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1045 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1004 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1015 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_15 VGND VPWR sky130_fd_sc_hd__fill_2
X_7247_ _7602_/Q la_data_in[96] _7247_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_49_26 VGND VPWR sky130_fd_sc_hd__decap_8
X_4459_ _4459_/A _4459_/B _4459_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_160_975 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_208 VGND VPWR sky130_fd_sc_hd__decap_12
X_7178_ _7604_/Q _7180_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_58_422 VGND VPWR sky130_fd_sc_hd__decap_12
X_6129_ _4320_/B _6128_/B _6101_/X _6129_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_46_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_959 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_1051 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_853 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_190 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1111 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_1189 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_823 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1136 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_806 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_385 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1106 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1109 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_86 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_867 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_147 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_232 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_883 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_511 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_724 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_663 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_50 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_482 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_107_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1235 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_806 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_485 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_349 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_236 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_820 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_127 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_330 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_864 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_80 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_464 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_867 VGND VPWR sky130_fd_sc_hd__decap_12
X_3830_ _4747_/A _3798_/B _3832_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_162_1239 VGND VPWR sky130_fd_sc_hd__decap_12
X_3761_ _3769_/A _3761_/B _3760_/Y _3761_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_13_580 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_861 VGND VPWR sky130_fd_sc_hd__decap_12
X_5500_ _5464_/X _5478_/X _5498_/X _5499_/X _5500_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_119_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_562 VGND VPWR sky130_fd_sc_hd__decap_12
X_6480_ wb_rst_i _6670_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_185_371 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_3692_ _4609_/A _4535_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_203_1269 VGND VPWR sky130_fd_sc_hd__decap_8
X_5431_ _5431_/A _5430_/X _5431_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_199_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_950 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1242 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_706 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_257 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_279 VGND VPWR sky130_fd_sc_hd__decap_12
X_5362_ _4695_/A _4505_/B _5363_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_142_920 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_227 VGND VPWR sky130_fd_sc_hd__decap_12
X_7101_ _6052_/A _7128_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_126_493 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_110 VGND VPWR sky130_fd_sc_hd__decap_12
X_4313_ _4256_/X _4307_/X _4311_/Y _4312_/X _4313_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_82_1218 VGND VPWR sky130_fd_sc_hd__decap_12
X_5293_ _5122_/X _5126_/X _5125_/X _5293_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_114_666 VGND VPWR sky130_fd_sc_hd__fill_2
X_7032_ _6967_/A la_data_in[64] _7032_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_102_828 VGND VPWR sky130_fd_sc_hd__decap_8
X_4244_ _4215_/X _4232_/X _4233_/X _4243_/X _4244_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_68_753 VGND VPWR sky130_fd_sc_hd__decap_8
X_4175_ _4172_/X _4174_/B _4174_/X _4175_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_95_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1076 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_583 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_959 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_406 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_812 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1103 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_288 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_806 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_322 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6816_ _6913_/A _6912_/A VGND VPWR sky130_fd_sc_hd__buf_1
XPHY_2129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7796_ _7796_/D _7796_/Q _7801_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_135 VGND VPWR sky130_fd_sc_hd__decap_12
X_6747_ _6747_/A _6747_/B _6747_/X VGND VPWR sky130_fd_sc_hd__and2_4
XPHY_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_850 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_809 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_27 VGND VPWR sky130_fd_sc_hd__decap_12
X_3959_ _3947_/Y _3958_/B _3959_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_211_478 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1112 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1006 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_883 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_574 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1066 VGND VPWR sky130_fd_sc_hd__fill_2
X_6678_ _6657_/X _6676_/X _6677_/Y _6678_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_17_1197 VGND VPWR sky130_fd_sc_hd__decap_12
X_5629_ _5614_/X _5620_/X _5627_/X _5628_/X _5629_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_191_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_577 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_739 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_994 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_611 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_430 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_761 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_625 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_1230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1121 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_753 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_1203 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_894 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_734 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_447 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_907 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_239 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_417 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_672 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_823 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_300 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_452 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_50 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_867 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_72 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_83 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_434 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_94 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_496 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_815 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_366 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_995 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_697 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_837 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1122 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_703 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_714 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_419 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1081 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_826 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1049 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_1224 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_76 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_959 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_425 VGND VPWR sky130_fd_sc_hd__fill_2
X_5980_ _5953_/X _5979_/X _5980_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_18_661 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_1000 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_597 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_288 VGND VPWR sky130_fd_sc_hd__decap_12
X_4931_ _4929_/X _4930_/X _4929_/X _4930_/X _4931_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_36_1006 VGND VPWR sky130_fd_sc_hd__fill_1
X_7650_ _7650_/D _6860_/A _7756_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_127_1123 VGND VPWR sky130_fd_sc_hd__decap_12
X_4862_ _5162_/A _4394_/B _4863_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_32_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_303 VGND VPWR sky130_fd_sc_hd__decap_12
X_6601_ la_data_in[30] _6601_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_75_1099 VGND VPWR sky130_fd_sc_hd__decap_12
X_3813_ _4645_/A _3813_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_177_135 VGND VPWR sky130_fd_sc_hd__decap_12
X_7581_ _7581_/HI la_data_out[108] VGND VPWR sky130_fd_sc_hd__conb_1
XANTENNA_15 _7276_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_4793_ _4793_/A _4793_/B _4793_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_162_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1011 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_703 VGND VPWR sky130_fd_sc_hd__decap_12
X_6532_ la_data_in[1] _6532_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_192_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_3744_ _7813_/Q _4613_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_118_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_381 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_544 VGND VPWR sky130_fd_sc_hd__decap_12
X_6463_ _6438_/X _6461_/X _6462_/Y _6463_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_203_1099 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_886 VGND VPWR sky130_fd_sc_hd__decap_8
X_5414_ _5347_/X _5351_/X _5347_/X _5351_/X _5414_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_173_374 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_739 VGND VPWR sky130_fd_sc_hd__decap_12
X_6394_ _6394_/A _6396_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_5345_ _5340_/X _5344_/X _5340_/X _5344_/X _5345_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_115_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_923 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_837 VGND VPWR sky130_fd_sc_hd__decap_12
X_5276_ _3773_/X _5275_/X _5276_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_99_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_293 VGND VPWR sky130_fd_sc_hd__decap_12
X_7015_ _6977_/X _7013_/X _7014_/Y _7015_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_101_135 VGND VPWR sky130_fd_sc_hd__decap_12
X_4227_ _4226_/A _4225_/X _4240_/A _4227_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_130_978 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_701 VGND VPWR sky130_fd_sc_hd__fill_1
X_4158_ _4118_/X _4119_/X _4118_/X _4119_/X _4158_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_56_734 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_210_1048 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_391 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_447 VGND VPWR sky130_fd_sc_hd__decap_8
X_4089_ _4072_/X _4088_/X _4072_/X _4088_/X _4089_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_83_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_417 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1182 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_44 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_642 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_664 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1245 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_995 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_242 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_1218 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7779_ _7779_/D _7779_/Q _7810_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_23_196 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_566 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_257 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1065 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_856 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_452 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_1173 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1014 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1088 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_288 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_480 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_236 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_93 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_450 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_293 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_105 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_820 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_511 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_190_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_1053 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1121 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_863 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_300 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_845 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_878 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_709 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_80 VGND VPWR sky130_fd_sc_hd__decap_12
X_5130_ _5130_/A _4903_/B _5130_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_97_623 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_645 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_293 VGND VPWR sky130_fd_sc_hd__decap_12
X_5061_ _5057_/X _5058_/X _5059_/Y _5060_/X _5061_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_97_678 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_818 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_870 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_317 VGND VPWR sky130_fd_sc_hd__decap_12
X_4012_ _4010_/X _4011_/X _4009_/X _4012_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_133_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_734 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_361 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_428 VGND VPWR sky130_fd_sc_hd__decap_12
X_5963_ _5963_/A _5963_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_203_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_581 VGND VPWR sky130_fd_sc_hd__decap_12
X_4914_ _4852_/X _4858_/X _4857_/X _4914_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_7702_ _6588_/X _7702_/Q _7696_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_209_1242 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_1253 VGND VPWR sky130_fd_sc_hd__decap_8
X_5894_ _5894_/A _5894_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_178_422 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_1275 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_444 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_623 VGND VPWR sky130_fd_sc_hd__decap_12
X_4845_ _4842_/X _4844_/X _4845_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7633_ _7100_/Y io_out[5] _7797_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_193_403 VGND VPWR sky130_fd_sc_hd__decap_12
X_7564_ _7564_/HI la_data_out[91] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_178_499 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_820 VGND VPWR sky130_fd_sc_hd__decap_8
X_4776_ _4847_/A _5123_/B _4779_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_53_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_166 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_105_1251 VGND VPWR sky130_fd_sc_hd__decap_12
X_6515_ _6515_/A _6515_/B _6515_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_158_190 VGND VPWR sky130_fd_sc_hd__decap_12
X_3727_ _4902_/A _4561_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_7495_ _7495_/HI la_data_out[22] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_162_801 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_683 VGND VPWR sky130_fd_sc_hd__decap_12
X_6446_ la_data_in[127] _6447_/B _6446_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_146_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_856 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_355 VGND VPWR sky130_fd_sc_hd__decap_8
X_6377_ wbs_dat_i[1] _6364_/B _6377_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_121_208 VGND VPWR sky130_fd_sc_hd__decap_12
X_5328_ _5298_/X _5327_/X _5298_/X _5327_/X _5328_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_115_794 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_422 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_1093 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_549 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_678 VGND VPWR sky130_fd_sc_hd__decap_12
X_5259_ _5099_/A _4778_/B _5259_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_75_306 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_1274 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_501 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_726 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_383 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_523 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_597 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_401 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_412 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_422 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1072 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_423 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_910 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_483 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1015 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_954 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1026 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_605 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_105 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_678 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_341 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_631 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_528 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1005 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_1182 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_1062 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_764 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_857 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_556 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1150 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_269 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_910 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_472 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_915 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_175_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_617 VGND VPWR sky130_fd_sc_hd__decap_12
X_4630_ _4624_/X _4629_/X _4628_/X _4630_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XPHY_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_1159 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_497 VGND VPWR sky130_fd_sc_hd__decap_12
X_4561_ _4561_/A _4479_/B _4561_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_6300_ _5977_/B _6300_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_7280_ _7256_/A _7280_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_155_171 VGND VPWR sky130_fd_sc_hd__decap_12
X_4492_ _4492_/A _4565_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_200_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_396 VGND VPWR sky130_fd_sc_hd__fill_1
X_6231_ _6229_/Y _6231_/B _7765_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_170_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1252 VGND VPWR sky130_fd_sc_hd__decap_12
X_6162_ _6147_/Y _6154_/Y _6162_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_170_1113 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_442 VGND VPWR sky130_fd_sc_hd__decap_12
X_5113_ _5108_/X _5112_/X _5111_/X _5113_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_112_764 VGND VPWR sky130_fd_sc_hd__decap_12
X_6093_ _3913_/Y _6091_/X _6092_/X _6093_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_57_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1119 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_1179 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_1110 VGND VPWR sky130_fd_sc_hd__decap_6
X_5044_ _4977_/X _4978_/X _4946_/X _4979_/X _5045_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_111_296 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_873 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_350 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_737 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1210 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6995_ _7647_/Q la_data_in[77] _6931_/X _6995_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_0_1265 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_1212 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1276 VGND VPWR sky130_fd_sc_hd__fill_1
X_5946_ _5946_/A _5945_/X _5946_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_90_1103 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_921 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_1245 VGND VPWR sky130_fd_sc_hd__decap_12
X_5877_ _5869_/X _5876_/X _5869_/X _5876_/X _5878_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_159_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_606 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_178_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_4828_ _3728_/X _4906_/B _4828_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7616_ _7210_/X _7616_/Q _7729_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4759_ _4759_/A _4758_/X _4759_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7547_ _7547_/HI la_data_out[74] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_181_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_525 VGND VPWR sky130_fd_sc_hd__decap_12
X_7478_ _7478_/HI la_data_out[5] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_4_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1013 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_32 VGND VPWR sky130_fd_sc_hd__decap_12
X_6429_ _6429_/A _6429_/B _6429_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_136_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_995 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_837 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_943 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_818 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_368 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1093 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_1172 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_895 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1018 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_827 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_394 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_337 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_220 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_242 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_762 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_286 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_773 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_297 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_83 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1020 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_650 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_468 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1135 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_483 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_685 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_442 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_615 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_497 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_339 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_1160 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_1130 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_654 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_501 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_208_676 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_843 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_1207 VGND VPWR sky130_fd_sc_hd__decap_12
X_5800_ _5785_/X _5791_/X _5798_/X _5799_/X _5801_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_35_578 VGND VPWR sky130_fd_sc_hd__decap_6
X_6780_ _6768_/X _6778_/X _6779_/Y _6780_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_3992_ _3966_/B _3968_/X _3991_/X _3994_/A VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_211_819 VGND VPWR sky130_fd_sc_hd__decap_12
X_5731_ _5731_/A _4901_/A _5731_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_200_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_329 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_128_1081 VGND VPWR sky130_fd_sc_hd__decap_12
X_5662_ _5658_/X _5659_/X _5660_/X _5661_/X _5662_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_176_745 VGND VPWR sky130_fd_sc_hd__decap_12
X_4613_ _4613_/A _4613_/B _4615_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_7401_ _7400_/Y _7387_/A _7777_/Q _7257_/X wbs_dat_o[31] VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_15_1251 VGND VPWR sky130_fd_sc_hd__fill_1
X_5593_ _5591_/X _5592_/X _5593_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_191_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_661 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_428 VGND VPWR sky130_fd_sc_hd__decap_12
X_7332_ _7332_/A _7321_/B _7332_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_116_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1126 VGND VPWR sky130_fd_sc_hd__decap_8
X_4544_ _4528_/X _4537_/X _4542_/X _4543_/X _4544_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_144_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1227 VGND VPWR sky130_fd_sc_hd__fill_1
X_7263_ io_in[6] _7263_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4475_ _4475_/A _4475_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_132_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_388 VGND VPWR sky130_fd_sc_hd__decap_8
X_6214_ _6212_/Y _6213_/X _6214_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_171_483 VGND VPWR sky130_fd_sc_hd__decap_4
X_7194_ _7163_/Y _7165_/B _7165_/X _7193_/X _7194_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_143_196 VGND VPWR sky130_fd_sc_hd__decap_12
X_6145_ _4309_/A _6103_/X _6144_/X _6145_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_6076_ _6317_/C _6308_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_39_851 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_607 VGND VPWR sky130_fd_sc_hd__decap_3
X_5027_ _5020_/Y _5021_/X _5023_/X _5027_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_85_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_117 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_556 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_662 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1051 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_898 VGND VPWR sky130_fd_sc_hd__decap_12
X_6978_ _6947_/Y _6949_/B _6949_/X _6977_/X _6978_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_179_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_44 VGND VPWR sky130_fd_sc_hd__decap_12
X_5929_ _5898_/X _5899_/X _5900_/X _5929_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_107_1121 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_1004 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_146_1181 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1075 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_924 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_726 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_979 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_737 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_439 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_611 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_509 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_154 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_407 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_309 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_938 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_426 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_556 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_887 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_386 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_93 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_1104 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_609 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_789 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_173_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_491 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_642 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_471 VGND VPWR sky130_fd_sc_hd__decap_8
X_4260_ _4769_/A _4328_/B _4260_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_119_1036 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_158_1096 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1233 VGND VPWR sky130_fd_sc_hd__decap_12
X_4191_ _4187_/X _4190_/Y _4187_/X _4190_/Y _4191_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_140_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_905 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_456 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_963 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_670 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_117 VGND VPWR sky130_fd_sc_hd__decap_12
X_6901_ _6912_/A _6874_/X _6901_/C _6901_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_82_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_342 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_211_32 VGND VPWR sky130_fd_sc_hd__decap_12
X_6832_ la_data_in[58] _6832_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_165_1034 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_846 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_87 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_1078 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_306 VGND VPWR sky130_fd_sc_hd__decap_12
X_3975_ _3973_/X _3974_/X _3975_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_6763_ _6727_/Y _6728_/Y _6762_/X _6763_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_206_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_879 VGND VPWR sky130_fd_sc_hd__decap_12
X_5714_ _5712_/X _5713_/X _5712_/X _5713_/X _5714_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_176_520 VGND VPWR sky130_fd_sc_hd__decap_12
X_6694_ _6913_/A _6694_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_149_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_907 VGND VPWR sky130_fd_sc_hd__decap_8
X_5645_ _5466_/X _5470_/X _5466_/X _5470_/X _5645_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_164_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_288 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_439 VGND VPWR sky130_fd_sc_hd__fill_1
X_5576_ _5573_/A _5572_/X _5575_/X _5576_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_145_951 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_1160 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_163_269 VGND VPWR sky130_fd_sc_hd__decap_12
X_4527_ _4474_/X _4510_/X _4474_/X _4510_/X _4527_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7315_ _7315_/A _7292_/B _7315_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_176_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1182 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_408 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_943 VGND VPWR sky130_fd_sc_hd__decap_3
X_4458_ _4452_/X _4457_/X _4456_/X _4458_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_7246_ _7238_/A _7246_/B _7245_/Y _7246_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_172_1027 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_678 VGND VPWR sky130_fd_sc_hd__decap_12
X_7177_ _7175_/Y _7177_/B _7177_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_4389_ _4351_/X _4352_/X _4351_/X _4352_/X _4389_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6128_ _4320_/B _6128_/B _6128_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_100_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_15 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_564 VGND VPWR sky130_fd_sc_hd__fill_1
X_6059_ _6332_/A _6059_/B _6059_/C _6059_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_46_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1090 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_821 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_1063 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_4214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_623 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_971 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1148 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_857 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_829 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_98 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_879 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_367 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_378 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_840 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_159 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_564 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_776 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_1181 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_556 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_642 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1211 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_910 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_280 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_954 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_1247 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_964 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_975 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_986 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1013 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_497 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_71 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1046 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_496 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1068 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_248 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_426 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_437 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1007 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_1067 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_922 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_459 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_876 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_109 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_898 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_4770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1259 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_520 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1081 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_518 VGND VPWR sky130_fd_sc_hd__fill_1
X_3760_ wbs_dat_i[18] _3790_/B _3760_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_13_592 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_873 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_406 VGND VPWR sky130_fd_sc_hd__fill_1
X_3691_ _4898_/A _4609_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_173_501 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_597 VGND VPWR sky130_fd_sc_hd__fill_1
X_5430_ _5099_/A _4492_/A _5430_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_69_1008 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_1019 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1038 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_962 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_578 VGND VPWR sky130_fd_sc_hd__fill_1
X_5361_ _4455_/A _4299_/X _5363_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_12_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_932 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_483 VGND VPWR sky130_fd_sc_hd__decap_3
X_4312_ _4256_/X _4307_/X _4256_/X _4307_/X _4312_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7100_ _7404_/A _7100_/B _7099_/X _7100_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_160_239 VGND VPWR sky130_fd_sc_hd__decap_12
X_5292_ _5292_/A _5292_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_141_453 VGND VPWR sky130_fd_sc_hd__decap_8
X_7031_ _7012_/A _6969_/X _7030_/Y _7031_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_206_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_367 VGND VPWR sky130_fd_sc_hd__decap_12
X_4243_ _4239_/X _4242_/X _4239_/X _4242_/X _4243_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_101_306 VGND VPWR sky130_fd_sc_hd__decap_12
X_4174_ _4172_/X _4174_/B _4174_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_136_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_562 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_618 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_1088 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_595 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_971 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_109 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1115 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6815_ _6795_/A _6815_/B _6814_/Y _6815_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_7795_ _7795_/D _7795_/Q _7797_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_211_435 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_367 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_91_1050 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6746_ la_data_in[34] _6747_/B VGND VPWR sky130_fd_sc_hd__inv_8
X_3958_ _3947_/Y _3958_/B _3958_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_195_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1124 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_1018 VGND VPWR sky130_fd_sc_hd__decap_12
X_3889_ _5198_/A _3897_/B _3891_/B VGND VPWR sky130_fd_sc_hd__and2_4
X_6677_ _6657_/X _6676_/X _6670_/X _6677_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_167_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_895 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_821 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_394 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_843 VGND VPWR sky130_fd_sc_hd__fill_1
X_5628_ _5614_/X _5620_/X _5614_/X _5620_/X _5628_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_191_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_589 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_898 VGND VPWR sky130_fd_sc_hd__decap_12
X_5559_ _5552_/X _5553_/X _5552_/X _5553_/X _5559_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_145_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_32 VGND VPWR sky130_fd_sc_hd__decap_12
X_7229_ _7193_/X _7228_/X _7212_/X _7229_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_104_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1250 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_637 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_1141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1242 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_708 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1248 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_746 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_459 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_919 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_651 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1_0_wb_clk_i clkbuf_2_0_1_wb_clk_i/X clkbuf_4_3_0_wb_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_3310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_684 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_835 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_312 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_40 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_51 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_199_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1073 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_51 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_62 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_73 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_879 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_84 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_446 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_378 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_175 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_350 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_540 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_726 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_551 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_940 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_450 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_239 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_1180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_194_1060 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_750 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_838 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1099 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_11 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_220 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_1236 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_532 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_565 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_971 VGND VPWR sky130_fd_sc_hd__decap_12
X_4930_ _4860_/X _4864_/X _4863_/X _4930_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_75_1012 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_993 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_963 VGND VPWR sky130_fd_sc_hd__decap_12
X_4861_ _5095_/A _4647_/B _4861_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_178_626 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_1135 VGND VPWR sky130_fd_sc_hd__decap_12
X_6600_ _6600_/A _6600_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_3812_ _4590_/A _4645_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_20_315 VGND VPWR sky130_fd_sc_hd__decap_12
X_4792_ _4780_/X _4782_/X _4779_/X _4792_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_7580_ _7580_/HI la_data_out[107] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_177_147 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_16 _7270_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_337 VGND VPWR sky130_fd_sc_hd__decap_12
X_3743_ _3743_/A _3769_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_6531_ _6531_/A _6531_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_119_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_832 VGND VPWR sky130_fd_sc_hd__decap_12
X_6462_ _6438_/X _6461_/X _6455_/X _6462_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_9_393 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_556 VGND VPWR sky130_fd_sc_hd__decap_4
X_5413_ _5408_/X _5412_/X _5411_/X _5413_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_6393_ _6391_/Y _6393_/B _6393_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_161_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1103 VGND VPWR sky130_fd_sc_hd__fill_1
X_5344_ _5343_/A _5343_/B _5343_/X _5344_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_173_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_1147 VGND VPWR sky130_fd_sc_hd__decap_12
X_5275_ _5533_/B _5275_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_130_935 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_849 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_1128 VGND VPWR sky130_fd_sc_hd__fill_1
X_4226_ _4226_/A _4225_/X _4240_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_7014_ _6977_/X _7013_/X _6999_/X _7014_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_101_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_916 VGND VPWR sky130_fd_sc_hd__decap_12
X_4157_ _4121_/X _4128_/X _4121_/X _4128_/X _4157_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_56_746 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_459 VGND VPWR sky130_fd_sc_hd__decap_12
X_4088_ _4073_/X _4079_/X _4080_/X _4087_/X _4088_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_209_590 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1112 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1243 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_56 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_924 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_1145 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1265 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_440 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_676 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_196_434 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_175 VGND VPWR sky130_fd_sc_hd__decap_8
X_7778_ _6146_/Y _4308_/A _7810_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6729_ _6727_/Y _6728_/Y _6727_/Y _6728_/Y _6794_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_137_512 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_383 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1028 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_868 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_558 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1217 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_497 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_318 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1185 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1067 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_1026 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_971 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_492 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_952 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_924 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_733 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_602 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_968 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_147 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_276 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_670 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1062 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_117 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1070 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_93 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1065 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_342 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_875 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_589 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_795 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_657 VGND VPWR sky130_fd_sc_hd__decap_12
X_5060_ _5057_/X _5058_/X _5057_/X _5058_/X _5060_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_42_1011 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_3 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_1191 VGND VPWR sky130_fd_sc_hd__decap_12
X_4011_ _4793_/A _4078_/B _4011_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_96_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_882 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_329 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_133_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_746 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_971 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_896 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_289 VGND VPWR sky130_fd_sc_hd__fill_1
X_5962_ _5955_/X _5961_/X _5963_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_7701_ _6591_/X _6525_/A _7707_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4913_ _4846_/X _4847_/X _4845_/X _4913_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_206_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_440 VGND VPWR sky130_fd_sc_hd__decap_12
X_5893_ _4741_/A _5443_/B _5893_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7632_ _7103_/X _7034_/A _7797_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4844_ _4844_/A _4844_/B _4844_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_178_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_415 VGND VPWR sky130_fd_sc_hd__decap_12
X_7563_ _7563_/HI la_data_out[90] VGND VPWR sky130_fd_sc_hd__conb_1
X_4775_ _5300_/B _5123_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_53_1184 VGND VPWR sky130_fd_sc_hd__decap_12
X_6514_ la_data_in[7] _6515_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_105_1263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1203 VGND VPWR sky130_fd_sc_hd__decap_12
X_3726_ _7815_/Q _4902_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_7494_ _7494_/HI la_data_out[21] VGND VPWR sky130_fd_sc_hd__conb_1
X_6445_ io_out[7] _6444_/X _6447_/B VGND VPWR sky130_fd_sc_hd__xnor2_4
XFILLER_49_1209 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_695 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_868 VGND VPWR sky130_fd_sc_hd__decap_12
X_6376_ _4782_/B _6345_/A _6378_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_161_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_924 VGND VPWR sky130_fd_sc_hd__fill_1
X_5327_ _5325_/X _5326_/X _5325_/X _5326_/X _5327_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_142_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_743 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_123 VGND VPWR sky130_fd_sc_hd__decap_12
X_5258_ _5253_/X _5257_/X _5256_/X _5258_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_57_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_871 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1250 VGND VPWR sky130_fd_sc_hd__decap_8
X_4209_ _4153_/X _4203_/X _4153_/X _4203_/X _4210_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_5189_ _5186_/X _5187_/X _5188_/X _5189_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_112_1223 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_351 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_395 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_535 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_1093 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_402 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1013 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_413 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_721 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_985 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1084 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_922 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_703 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_495 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_123 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_966 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_489 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_617 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_117 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_459 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_802 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_353 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_721 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_635 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_399 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_191_1074 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_657 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_819 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_605 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_1099 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_616 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_798 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_705 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_440 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1252 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1143 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1026 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_484 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_1274 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1116 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_292 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_629 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_32 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_487 VGND VPWR sky130_fd_sc_hd__fill_1
X_4560_ _4551_/X _4557_/X _4558_/X _4559_/X _4560_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_198_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_76 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_353 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_813 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_301 VGND VPWR sky130_fd_sc_hd__decap_4
X_4491_ _4491_/A _4492_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_183_470 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1059 VGND VPWR sky130_fd_sc_hd__decap_8
X_6230_ _5292_/Y _6117_/X _6190_/X _6231_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_143_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_1182 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_922 VGND VPWR sky130_fd_sc_hd__decap_8
X_6161_ _5032_/B _6153_/X _6161_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_48_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_220 VGND VPWR sky130_fd_sc_hd__decap_12
X_5112_ _5111_/A _5110_/X _5111_/X _5112_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_170_1125 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_808 VGND VPWR sky130_fd_sc_hd__decap_12
X_6092_ _6068_/A _6092_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_454 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_318 VGND VPWR sky130_fd_sc_hd__decap_12
X_5043_ _5035_/X _5036_/X _5035_/X _5036_/X _5045_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_362 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_168_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1222 VGND VPWR sky130_fd_sc_hd__decap_12
X_6994_ _6923_/A _6994_/B _6994_/C _7648_/D VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_81_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_708 VGND VPWR sky130_fd_sc_hd__decap_12
X_5945_ _7796_/Q _7730_/Q _5945_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_179_721 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_1262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1115 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_398 VGND VPWR sky130_fd_sc_hd__decap_12
X_5876_ _5874_/X _5875_/X _5874_/X _5875_/X _5876_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_167_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1254 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1276 VGND VPWR sky130_fd_sc_hd__fill_1
X_7615_ _7214_/X _7615_/Q _7729_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_166_415 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_139_629 VGND VPWR sky130_fd_sc_hd__decap_12
X_4827_ _4612_/B _4906_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_138_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_908 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_245 VGND VPWR sky130_fd_sc_hd__decap_12
X_7546_ _7546_/HI la_data_out[73] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_105_1060 VGND VPWR sky130_fd_sc_hd__decap_8
X_4758_ _4547_/A _4758_/B _4758_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_147_684 VGND VPWR sky130_fd_sc_hd__decap_6
X_3709_ _6038_/A _6038_/B _3709_/C _3709_/D _6323_/A VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_88_1044 VGND VPWR sky130_fd_sc_hd__decap_12
X_7477_ _7477_/HI la_data_out[4] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_175_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_4689_ _4676_/X _4686_/X _4687_/X _4688_/X _4689_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_179_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1025 VGND VPWR sky130_fd_sc_hd__decap_12
X_6428_ _6415_/Y _6417_/B _6417_/X _6427_/X _6429_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_135_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_410 VGND VPWR sky130_fd_sc_hd__decap_12
X_6359_ _4293_/X _6373_/B _6361_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_0_314 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_955 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1217 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1111 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1020 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_811 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_806 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_204 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_839 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_74 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_877 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_349 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_210 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_220 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_232 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_410 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_243 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_713 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_265 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_938 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_977 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_276 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_287 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_298 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_785 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_448 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_95 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_790 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_529 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_581 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_697 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_540 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_454 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_121_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1153 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1219 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_80 VGND VPWR sky130_fd_sc_hd__decap_12
X_3991_ _3991_/A _3990_/X _3991_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_90_685 VGND VPWR sky130_fd_sc_hd__decap_12
X_5730_ _4743_/A _4363_/A _5730_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_16_793 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_905 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1093 VGND VPWR sky130_fd_sc_hd__decap_12
X_5661_ _5649_/X _5650_/X _5649_/X _5650_/X _5661_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_176_757 VGND VPWR sky130_fd_sc_hd__decap_6
X_7400_ io_in[37] _7400_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4612_ _4612_/A _4612_/B _4612_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_175_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1025 VGND VPWR sky130_fd_sc_hd__decap_8
X_5592_ _5200_/A _4145_/A _5592_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_191_727 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_141_1271 VGND VPWR sky130_fd_sc_hd__decap_6
X_7331_ _5639_/A _7309_/X _7327_/X _7330_/Y wbs_dat_o[11] VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_190_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_684 VGND VPWR sky130_fd_sc_hd__decap_12
X_4543_ _4528_/X _4537_/X _4528_/X _4537_/X _4543_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_144_621 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_654 VGND VPWR sky130_fd_sc_hd__decap_8
X_7262_ _7370_/A _7262_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_117_879 VGND VPWR sky130_fd_sc_hd__decap_12
X_4474_ _4458_/X _4464_/X _4472_/X _4473_/X _4474_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_209_98 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_304 VGND VPWR sky130_fd_sc_hd__fill_1
X_6213_ _5582_/X _6199_/X _5581_/A _6213_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_132_849 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_326 VGND VPWR sky130_fd_sc_hd__fill_1
X_7193_ _7166_/Y _7168_/B _7168_/X _7192_/X _7193_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_98_741 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1020 VGND VPWR sky130_fd_sc_hd__decap_12
X_6144_ _6144_/A _6144_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_58_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_785 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_402 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_936 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_947 VGND VPWR sky130_fd_sc_hd__fill_1
X_6075_ _6185_/A _6074_/X _6075_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_5026_ _5018_/X _5019_/X _5024_/X _5025_/X _5026_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_22_1234 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_619 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_129 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_28 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_827 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_568 VGND VPWR sky130_fd_sc_hd__decap_12
X_6977_ _6952_/A _6952_/B _6952_/X _6976_/X _6977_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XPHY_3739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_337 VGND VPWR sky130_fd_sc_hd__decap_12
X_5928_ _5923_/X _5924_/X _5923_/X _5924_/X _5928_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_702 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_179_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_831 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_426 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_5859_ _5824_/X _5840_/X _5841_/X _5859_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_55_1087 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1008 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_936 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1177 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_971 VGND VPWR sky130_fd_sc_hd__decap_12
X_7529_ _7529_/HI la_data_out[56] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_5_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_805 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_613 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_337 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_679 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_1206 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1036 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_419 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_917 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_608 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_899 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_516 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_696 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_398 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1154 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_201_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_521 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_1127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_251 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_745 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_576 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_971 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_173_727 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_200_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_337 VGND VPWR sky130_fd_sc_hd__decap_12
X_4190_ _4190_/A _4189_/X _4190_/Y VGND VPWR sky130_fd_sc_hd__xnor2_4
XFILLER_68_914 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_1245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_1204 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_402 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_882 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_936 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1248 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_811 VGND VPWR sky130_fd_sc_hd__decap_12
X_6900_ _6874_/A _6873_/X _6901_/C VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_209_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_682 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1021 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_169_1160 VGND VPWR sky130_fd_sc_hd__decap_12
X_6831_ _7660_/Q _6833_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_211_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_685 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_899 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1008 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1221 VGND VPWR sky130_fd_sc_hd__decap_12
X_6762_ _6794_/A _6761_/X _6762_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_3974_ _4612_/A _4218_/B _3974_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_210_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_702 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1032 VGND VPWR sky130_fd_sc_hd__decap_12
X_5713_ _5639_/Y _5640_/X _5639_/Y _5640_/X _5713_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6693_ _6052_/A _6913_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_176_532 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1238 VGND VPWR sky130_fd_sc_hd__decap_12
X_5644_ _5633_/X _5634_/X _5632_/Y _5635_/X _5644_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_164_727 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_513 VGND VPWR sky130_fd_sc_hd__decap_12
X_5575_ _5573_/Y _5574_/Y _5575_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_7314_ _5807_/A _7309_/X _7310_/X _7313_/Y wbs_dat_o[8] VGND VPWR sky130_fd_sc_hd__a211o_4
Xclkbuf_4_3_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/A _7754_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_4526_ _4511_/X _4517_/X _4524_/X _4525_/X _4526_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_105_805 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_1142 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_676 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_1194 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_911 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1036 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_304 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_1115 VGND VPWR sky130_fd_sc_hd__decap_12
X_7245_ _7245_/A _7184_/X _7245_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_4457_ _4456_/A _4456_/B _4456_/X _4457_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_171_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_495 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1039 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_903 VGND VPWR sky130_fd_sc_hd__decap_12
X_7176_ la_data_in[99] _7177_/B VGND VPWR sky130_fd_sc_hd__inv_8
X_4388_ _4373_/X _4374_/X _4373_/X _4374_/X _4388_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_59_936 VGND VPWR sky130_fd_sc_hd__fill_1
X_6127_ _6123_/Y _6133_/B _4447_/B _6128_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_100_532 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1020 VGND VPWR sky130_fd_sc_hd__decap_8
X_6058_ _3909_/Y _6058_/B _6059_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_65_38 VGND VPWR sky130_fd_sc_hd__decap_12
X_5009_ _4992_/X _5008_/X _4992_/X _5008_/X _5009_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_27_833 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_4204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_855 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_983 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_825 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_162 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_606 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_184 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_398 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_59 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_521 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_59 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_571 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_852 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_407 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_576 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1160 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_440 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_760 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_269 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_1207 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_977 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_431 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_679 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_442 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_453 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_464 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_475 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1025 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_83 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_703 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_800 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_833 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_449 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_1175 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_934 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_685 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_335 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_177_318 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1060 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_198_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_672 VGND VPWR sky130_fd_sc_hd__decap_12
X_3690_ _4820_/A _4898_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_146_727 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_524 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_790 VGND VPWR sky130_fd_sc_hd__decap_3
X_5360_ _4747_/A _4366_/B _5360_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_127_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_771 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_4311_ _4308_/A _4304_/Y _4310_/X _4311_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_5_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_944 VGND VPWR sky130_fd_sc_hd__fill_2
X_5291_ _5136_/X _5151_/X _5121_/X _5152_/X _5291_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_153_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_123 VGND VPWR sky130_fd_sc_hd__decap_12
X_7030_ _7030_/A _6968_/X _7030_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_4242_ _4240_/X _4241_/X _4240_/X _4241_/X _4242_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_142_988 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_379 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_733 VGND VPWR sky130_fd_sc_hd__fill_1
X_4173_ _4494_/A _4923_/B _4174_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_67_210 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_917 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_405 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_758 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_983 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_825 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6814_ _6814_/A _6814_/B _6814_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XPHY_2109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_121 VGND VPWR sky130_fd_sc_hd__decap_8
X_7794_ _7794_/D _6319_/A _7746_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_196_616 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_447 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_154 VGND VPWR sky130_fd_sc_hd__decap_12
X_6745_ _6745_/A _6747_/A VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3957_ _3957_/A _3956_/X _3958_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_143_1141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_198 VGND VPWR sky130_fd_sc_hd__decap_12
X_6676_ _6609_/A la_data_in[27] _6611_/X _6676_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_137_716 VGND VPWR sky130_fd_sc_hd__fill_1
X_3888_ _5233_/A _5198_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_176_362 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_5627_ _5624_/X _5625_/X _5626_/X _5627_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_178_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_557 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_440 VGND VPWR sky130_fd_sc_hd__fill_1
X_5558_ _5554_/X _5557_/X _5554_/X _5557_/X _5558_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_105_602 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_624 VGND VPWR sky130_fd_sc_hd__decap_12
X_4509_ _4502_/X _4508_/X _4502_/X _4508_/X _4509_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_133_944 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_5489_ _5486_/X _5487_/X _5501_/A _5489_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_160_741 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_977 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_668 VGND VPWR sky130_fd_sc_hd__decap_3
X_7228_ _7609_/Q la_data_in[103] _7165_/X _7228_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_133_988 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_605 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_700 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_487 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1153 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_733 VGND VPWR sky130_fd_sc_hd__decap_12
X_7159_ _7157_/Y _7158_/Y _7157_/Y _7158_/Y _7224_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_101_830 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_1189 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_758 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_4012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_257 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_663 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_30 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_904 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_471 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_791 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_696 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_41 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_847 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_324 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_52 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_63 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_476 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_74 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1085 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_1036 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_346 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_85 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_74 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_96 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1203 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_362 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_513 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_1179 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_516 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_771 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_495 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_1045 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_251 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_261 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_272 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_349 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_283 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_294 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_1248 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_714 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_720 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_706 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_731 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_577 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_983 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_151 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1024 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_605 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_184 VGND VPWR sky130_fd_sc_hd__decap_12
X_4860_ _5099_/A _4653_/B _4860_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_75_1057 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_638 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_80 VGND VPWR sky130_fd_sc_hd__decap_12
X_3811_ _3811_/A _4590_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_32_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_830 VGND VPWR sky130_fd_sc_hd__decap_12
X_4791_ _4738_/X _4767_/X _4789_/X _4790_/X _4791_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_207_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_327 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_17 _7288_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_177_159 VGND VPWR sky130_fd_sc_hd__decap_12
X_6530_ _6530_/A _6530_/B _6530_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_3742_ _6144_/A _3743_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_174_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_727 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_158_373 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_6461_ _6394_/A la_data_in[122] _6396_/X _6461_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_174_844 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1090 VGND VPWR sky130_fd_sc_hd__decap_8
X_5412_ _5409_/X _5410_/X _5411_/X _5412_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_6392_ la_data_in[123] _6393_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_127_771 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_410 VGND VPWR sky130_fd_sc_hd__decap_12
X_5343_ _5343_/A _5343_/B _5343_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_99_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1265 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_605 VGND VPWR sky130_fd_sc_hd__decap_8
X_5274_ _5261_/X _5274_/B _5274_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_7013_ _6947_/A la_data_in[71] _6949_/X _7013_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_4225_ _4519_/A _4591_/B _4225_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_101_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_928 VGND VPWR sky130_fd_sc_hd__decap_12
X_4156_ _4130_/X _4140_/X _4130_/X _4140_/X _4156_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_660 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_427 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_758 VGND VPWR sky130_fd_sc_hd__decap_4
X_4087_ _4086_/A _4085_/X _4086_/X _4087_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_55_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1124 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_68 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1157 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_211 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_7777_ _7777_/D _7777_/Q _7774_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1269 VGND VPWR sky130_fd_sc_hd__decap_8
X_4989_ _4986_/A _4985_/X _4988_/Y _4989_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XPHY_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6728_ la_data_in[40] _6728_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_524 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_395 VGND VPWR sky130_fd_sc_hd__decap_12
X_6659_ _6606_/Y _6608_/B _6608_/X _6658_/X _6659_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_165_855 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1120 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1062 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1270 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_728 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_983 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_780 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_611 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_936 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_964 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_745 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_947 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_154 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_997 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_614 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_187 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_468 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_669 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_682 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1074 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1082 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_129 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1044 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_894 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_877 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_505 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_887 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_741 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_327 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_1061 VGND VPWR sky130_fd_sc_hd__decap_12
X_4010_ _4007_/X _4008_/X _4009_/X _4010_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_77_371 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1203 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_758 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_577 VGND VPWR sky130_fd_sc_hd__decap_12
X_5961_ _5956_/Y _5958_/X _5959_/X _5960_/X _5961_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_18_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_931 VGND VPWR sky130_fd_sc_hd__decap_12
X_7700_ _7700_/D _7700_/Q _7707_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_179_903 VGND VPWR sky130_fd_sc_hd__decap_12
X_4912_ _4893_/X _4911_/X _4893_/X _4911_/X _4912_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_5892_ _5890_/X _5891_/X _5889_/X _5892_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_80_569 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_452 VGND VPWR sky130_fd_sc_hd__decap_6
X_7631_ _7631_/D _7037_/A _7729_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4843_ _4843_/A _4844_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_61_794 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_485 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_647 VGND VPWR sky130_fd_sc_hd__decap_12
X_7562_ _7562_/HI la_data_out[89] VGND VPWR sky130_fd_sc_hd__conb_1
X_4774_ _4769_/X _4773_/X _4772_/X _4774_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_119_502 VGND VPWR sky130_fd_sc_hd__decap_12
X_6513_ _7705_/Q _6515_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_3725_ _3733_/A _3725_/B _3724_/Y _3725_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_53_1196 VGND VPWR sky130_fd_sc_hd__decap_12
X_7493_ _7493_/HI la_data_out[20] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_119_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_1275 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_1106 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1215 VGND VPWR sky130_fd_sc_hd__decap_12
X_6444_ _6382_/Y _6383_/Y _6450_/B _6444_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_175_1207 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_398 VGND VPWR sky130_fd_sc_hd__decap_12
X_6375_ _6381_/A _6375_/B _6374_/Y _7732_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_115_741 VGND VPWR sky130_fd_sc_hd__fill_1
X_5326_ _5195_/X _5209_/X _5153_/X _5210_/X _5326_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_161_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1062 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_785 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_593 VGND VPWR sky130_fd_sc_hd__decap_12
X_5257_ _5254_/X _5255_/X _5256_/X _5257_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_87_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_1123 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_4208_ _4200_/X _4201_/X _4202_/X _4208_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_5188_ _5186_/X _5187_/X _5188_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_112_1235 VGND VPWR sky130_fd_sc_hd__decap_12
X_4139_ _3914_/A _4143_/A _4179_/A _4139_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_83_341 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_769 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_875 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_363 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_920 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_189_27 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_403 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_569 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1011 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_441 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_414 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_1025 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1082 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_733 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1096 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_934 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1047 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_715 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_185_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_658 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_135 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1203 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_145_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_629 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_129 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_64 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_857 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1192 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1023 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1031 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_3_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1004 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_733 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_628 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_837 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_801 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_566 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_257 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_717 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_931 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1016 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_1155 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1128 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1188 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_44 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_855 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_680 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_674 VGND VPWR sky130_fd_sc_hd__decap_3
X_4490_ _5835_/B _4491_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_171_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_482 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_7_684 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_346 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_154 VGND VPWR sky130_fd_sc_hd__decap_12
X_6160_ _6156_/X _6157_/Y _6159_/X _7777_/D VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_40_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_880 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_174_1262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1276 VGND VPWR sky130_fd_sc_hd__fill_1
X_5111_ _5111_/A _5110_/X _5111_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_98_956 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_135 VGND VPWR sky130_fd_sc_hd__decap_12
X_6091_ _6158_/A _6091_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_111_232 VGND VPWR sky130_fd_sc_hd__decap_12
X_5042_ _5039_/A _5040_/A _5041_/X _5042_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_112_788 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_265 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_661 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_672 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_300 VGND VPWR sky130_fd_sc_hd__decap_12
X_6993_ _6993_/A _6986_/X _6994_/C VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_19_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1234 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_867 VGND VPWR sky130_fd_sc_hd__decap_12
X_5944_ _5935_/Y _5936_/X _5935_/Y _5936_/X _5944_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_1252 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_569 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1041 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_179_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1052 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1274 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_1233 VGND VPWR sky130_fd_sc_hd__decap_4
X_5875_ _5845_/Y _5846_/X _5845_/Y _5846_/X _5875_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_1127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_293 VGND VPWR sky130_fd_sc_hd__decap_12
X_4826_ _4823_/X _4824_/X _4825_/X _4826_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_7614_ _7217_/X _7614_/Q _7785_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_178_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_427 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_7545_ _7545_/HI la_data_out[72] VGND VPWR sky130_fd_sc_hd__conb_1
X_4757_ _4590_/A _4757_/B _4759_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_147_641 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_257 VGND VPWR sky130_fd_sc_hd__decap_12
X_3708_ wbs_adr_i[4] _3700_/X _3707_/X _3709_/D VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_119_365 VGND VPWR sky130_fd_sc_hd__fill_1
X_7476_ _7476_/HI la_data_out[3] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_174_471 VGND VPWR sky130_fd_sc_hd__fill_1
X_4688_ _4676_/X _4686_/X _4676_/X _4686_/X _4688_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_88_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_110 VGND VPWR sky130_fd_sc_hd__decap_12
X_6427_ _6418_/Y _6420_/B _6420_/X _6426_/X _6427_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_179_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_912 VGND VPWR sky130_fd_sc_hd__decap_3
X_6358_ _6340_/A _6373_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_68_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_304 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_733 VGND VPWR sky130_fd_sc_hd__decap_12
X_5309_ _5307_/X _5308_/X _5307_/X _5308_/X _5309_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_89_967 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_191_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_6289_ _5984_/Y _6288_/X _6289_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_89_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_563 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_566 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_508 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_322 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_867 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_200 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_208 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_211 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_794 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_233 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_422 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_255 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_916 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_277 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_725 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_989 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_288 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_299 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_556 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_758 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_630 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_437 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1150 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_1082 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1172 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_335 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_964 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_806 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_560 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_153 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_477 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1165 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_689 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1198 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_867 VGND VPWR sky130_fd_sc_hd__decap_6
X_3990_ _3984_/X _3987_/X _3988_/Y _3989_/X _3990_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_206_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_697 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_219 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_742 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_928 VGND VPWR sky130_fd_sc_hd__decap_12
X_5660_ _5658_/X _5659_/X _5658_/X _5659_/X _5660_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_200_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_80 VGND VPWR sky130_fd_sc_hd__decap_12
X_4611_ _4608_/X _4609_/X _4813_/B _4611_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_30_274 VGND VPWR sky130_fd_sc_hd__fill_1
X_5591_ _5341_/A _4277_/A _5591_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_157_961 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_11 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1264 VGND VPWR sky130_fd_sc_hd__decap_12
X_7330_ _3813_/X _7322_/X _7329_/X _7330_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
X_4542_ _4538_/X _4539_/X _4540_/Y _4541_/X _4542_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_8_971 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_696 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_633 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_110 VGND VPWR sky130_fd_sc_hd__decap_12
X_7261_ _7261_/A _7370_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_85_1218 VGND VPWR sky130_fd_sc_hd__fill_2
X_4473_ _4458_/X _4464_/X _4458_/X _4464_/X _4473_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6212_ _5576_/X _6212_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_89_208 VGND VPWR sky130_fd_sc_hd__decap_12
X_7192_ _7169_/Y _7170_/Y _7236_/B _7192_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_125_891 VGND VPWR sky130_fd_sc_hd__decap_4
X_6143_ _6024_/Y _4451_/X _6024_/Y _4451_/X _6143_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_174_1081 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_135_1032 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_703 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_883 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_797 VGND VPWR sky130_fd_sc_hd__decap_8
X_6074_ _6256_/B _6061_/X _6072_/Y _3911_/Y _6073_/X _6074_/X VGND VPWR sky130_fd_sc_hd__o32a_4
X_5025_ _5018_/X _5019_/X _5018_/X _5019_/X _5025_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_22_1246 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_823 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_480 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_806 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_3707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1031 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_839 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_141 VGND VPWR sky130_fd_sc_hd__decap_12
X_6976_ _6953_/Y _6954_/Y _6975_/X _6976_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_13_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1086 VGND VPWR sky130_fd_sc_hd__decap_12
X_5927_ _5910_/X _5926_/X _5985_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_94_1093 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_1052 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_574 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_68 VGND VPWR sky130_fd_sc_hd__decap_12
X_5858_ _5853_/X _5854_/X _5853_/X _5854_/X _5858_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_166_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_854 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1156 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_1099 VGND VPWR sky130_fd_sc_hd__decap_12
X_4809_ _4579_/X _4585_/X _4545_/X _4586_/X _4809_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_194_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1069 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_1189 VGND VPWR sky130_fd_sc_hd__decap_12
X_5789_ _5789_/A _5789_/B _5789_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_10_959 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_898 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_983 VGND VPWR sky130_fd_sc_hd__decap_12
X_7528_ _7528_/HI la_data_out[55] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_135_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_7459_ _7459_/HI io_out[24] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_134_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1113 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_658 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_1181 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_156 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1048 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_406 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_970 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_428 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_672 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_311 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_525 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_193 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_867 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_205_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_883 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_257 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_1133 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_419 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_828 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1038 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_891 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1216 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_414 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_436 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_910 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_209_932 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_943 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_631 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1172 VGND VPWR sky130_fd_sc_hd__decap_8
X_6830_ _6830_/A _6830_/B _6830_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_211_56 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_697 VGND VPWR sky130_fd_sc_hd__decap_12
X_6761_ _6730_/Y _6732_/B _6732_/X _6760_/X _6761_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_3973_ _3728_/X _3950_/B _3973_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_91_1233 VGND VPWR sky130_fd_sc_hd__decap_12
X_5712_ _5700_/X _5701_/X _5695_/X _5702_/X _5712_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_210_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_714 VGND VPWR sky130_fd_sc_hd__decap_12
X_6692_ _6650_/X _6689_/X _6691_/Y _6692_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_206_1044 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_550 VGND VPWR sky130_fd_sc_hd__decap_12
X_5643_ _5631_/X _5636_/X _5641_/X _5642_/X _5643_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_149_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_577 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_164_739 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_117_600 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_1020 VGND VPWR sky130_fd_sc_hd__decap_12
X_5574_ _5572_/X _5574_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_191_525 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_611 VGND VPWR sky130_fd_sc_hd__decap_8
X_7313_ _5420_/A _7293_/X _7312_/X _7313_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
X_4525_ _4511_/X _4517_/X _4511_/X _4517_/X _4525_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_176_1121 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_154 VGND VPWR sky130_fd_sc_hd__decap_12
X_7244_ _7186_/X _7242_/X _7243_/Y _7244_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_160_923 VGND VPWR sky130_fd_sc_hd__decap_12
X_4456_ _4456_/A _4456_/B _4456_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_176_1165 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1127 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_349 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_131_135 VGND VPWR sky130_fd_sc_hd__decap_12
X_7175_ _7605_/Q _7175_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4387_ _4379_/X _4380_/X _4379_/X _4380_/X _4387_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_86_712 VGND VPWR sky130_fd_sc_hd__decap_8
X_6126_ _6125_/X _6133_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_86_767 VGND VPWR sky130_fd_sc_hd__decap_12
X_6057_ _6057_/A _6055_/X _6057_/C _6057_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_74_918 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1070 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_970 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_1262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_672 VGND VPWR sky130_fd_sc_hd__decap_3
X_5008_ _4993_/X _5002_/X _5006_/X _5007_/X _5008_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_113_1160 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_588 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_428 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_845 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_867 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_995 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_837 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_174 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_618 VGND VPWR sky130_fd_sc_hd__fill_1
X_6959_ _7637_/Q _6959_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_2825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_27 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_32 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_533 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_909 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_588 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_419 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_931 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_738 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_226 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_772 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_900 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_911 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1219 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_922 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1107 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_496 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_150_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_933 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_509 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_861 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1060 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_999 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_745 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_767 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_406 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1069 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1187 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_193 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_344 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1206 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_697 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_536 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_396 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_598 VGND VPWR sky130_fd_sc_hd__decap_12
X_4310_ _4309_/X _4310_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_5290_ _5068_/X _5069_/X _5062_/Y _5070_/X _5290_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_153_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_658 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_135 VGND VPWR sky130_fd_sc_hd__decap_12
X_4241_ _4180_/X _4185_/X _4180_/X _4185_/X _4241_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_84_1081 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_56 VGND VPWR sky130_fd_sc_hd__decap_12
X_4172_ _4168_/X _4170_/X _4171_/X _4172_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_171_1062 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_222 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_704 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_929 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_995 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_623 VGND VPWR sky130_fd_sc_hd__decap_12
X_6813_ _6753_/X _6809_/X _6812_/Y _6813_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_211_404 VGND VPWR sky130_fd_sc_hd__decap_12
X_7793_ _7793_/D _7348_/A _7785_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3956_ _3943_/X _3946_/Y _3947_/Y _3956_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_6744_ _6744_/A _6744_/B _6744_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_17_1123 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_459 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1191 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_188_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1153 VGND VPWR sky130_fd_sc_hd__decap_6
X_6675_ _6658_/X _6673_/X _6674_/Y _6675_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_3887_ _5178_/A _5233_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_31_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1069 VGND VPWR sky130_fd_sc_hd__fill_2
X_5626_ _5624_/X _5625_/X _5626_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_176_374 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_569 VGND VPWR sky130_fd_sc_hd__decap_8
X_5557_ _5555_/X _5556_/X _5555_/X _5556_/X _5557_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_3_708 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_208 VGND VPWR sky130_fd_sc_hd__decap_12
X_4508_ _4503_/X _4507_/X _4506_/X _4508_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_145_794 VGND VPWR sky130_fd_sc_hd__decap_8
X_5488_ _5486_/X _5487_/X _5501_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_132_422 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_636 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_956 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_753 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_444 VGND VPWR sky130_fd_sc_hd__decap_12
X_4439_ _4388_/X _4433_/X _4437_/X _4438_/X _4439_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_7227_ _7210_/A _7227_/B _7226_/Y _7227_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_160_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1252 VGND VPWR sky130_fd_sc_hd__decap_6
X_7158_ la_data_in[105] _7158_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_24_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_1274 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_745 VGND VPWR sky130_fd_sc_hd__decap_8
X_6109_ _6308_/B _6109_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_112_190 VGND VPWR sky130_fd_sc_hd__decap_12
X_7089_ _7117_/A _7088_/X _7118_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_58_255 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1228 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_597 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_480 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_962 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_910 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_20 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_612 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1042 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_42 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1004 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_100 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_53 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_64 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_75 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_358 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_86 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_105 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_97 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_86 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_459 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_892 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_520 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1275 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_168_886 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_993 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_502 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_525 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_74 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_157_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_901 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_783 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_1013 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_251 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_726 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_428 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1090 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_743 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_163 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1036 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_196 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_75_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3810_ _7805_/Q _3811_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_61_987 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_818 VGND VPWR sky130_fd_sc_hd__decap_12
X_4790_ _4738_/X _4767_/X _4738_/X _4767_/X _4790_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_32_166 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1003 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_18 _7295_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3741_ _3733_/A _3741_/B _3740_/Y _3741_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_13_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_340 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_812 VGND VPWR sky130_fd_sc_hd__decap_12
X_6460_ _6439_/X _6458_/X _6459_/Y _7725_/D VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_158_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_322 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_856 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1020 VGND VPWR sky130_fd_sc_hd__decap_12
X_5411_ _5409_/X _5410_/X _5411_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_51_1080 VGND VPWR sky130_fd_sc_hd__fill_1
X_6391_ _7725_/Q _6391_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_133_208 VGND VPWR sky130_fd_sc_hd__decap_12
X_5342_ _5233_/A _4854_/B _5343_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_127_794 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_114_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_1135 VGND VPWR sky130_fd_sc_hd__decap_12
X_5273_ _5230_/X _5251_/X _5271_/X _5272_/X _5273_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_142_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_306 VGND VPWR sky130_fd_sc_hd__decap_12
X_7012_ _7012_/A _7012_/B _7012_/C _7012_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_4224_ _4485_/A _4590_/B _4226_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_102_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_907 VGND VPWR sky130_fd_sc_hd__decap_8
X_4155_ _4142_/X _4148_/X _4142_/X _4148_/X _4155_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_110_650 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_715 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_512 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1221 VGND VPWR sky130_fd_sc_hd__decap_6
X_4086_ _4086_/A _4085_/X _4086_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_23_1160 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_450 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_239 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1215 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_689 VGND VPWR sky130_fd_sc_hd__decap_12
X_7776_ _7776_/D _4434_/A _7774_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_306 VGND VPWR sky130_fd_sc_hd__decap_12
X_4988_ _4987_/X _4988_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_609 VGND VPWR sky130_fd_sc_hd__fill_1
X_6727_ _6727_/A _6727_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_3939_ _4653_/B _4328_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_165_801 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_661 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_300 VGND VPWR sky130_fd_sc_hd__decap_12
X_6658_ _6611_/A _6611_/B _6611_/X _6657_/X _6658_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_137_536 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1024 VGND VPWR sky130_fd_sc_hd__fill_1
X_5609_ _5607_/X _5608_/X _5609_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_30_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_366 VGND VPWR sky130_fd_sc_hd__decap_12
X_6589_ _6525_/A la_data_in[3] _6527_/X _6589_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_3_516 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_720 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_328 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_531 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_851 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1074 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_759 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_545 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_932 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_792 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_757 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_166 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_626 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_199 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1170 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_840 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_300 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1094 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_884 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_361 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_321 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_855 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1146 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_517 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_697 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_899 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_764 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_306 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_583 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_339 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_593 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1073 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_501 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_383 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_269 VGND VPWR sky130_fd_sc_hd__decap_12
X_5960_ _5956_/Y _5958_/X _5956_/Y _5958_/X _5960_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_168_1248 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_589 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_483 VGND VPWR sky130_fd_sc_hd__decap_12
X_4911_ _4894_/X _4910_/X _4894_/X _4910_/X _4911_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_52_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_943 VGND VPWR sky130_fd_sc_hd__decap_3
X_5891_ _3877_/A _5835_/B _5891_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7630_ _7630_/D _7040_/A _7729_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_209_1267 VGND VPWR sky130_fd_sc_hd__decap_8
X_4842_ _3763_/A _4915_/B _4842_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4773_ _4772_/A _4771_/X _4772_/X _4773_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_7561_ _7561_/HI la_data_out[88] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_92_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_514 VGND VPWR sky130_fd_sc_hd__decap_12
X_3724_ wbs_dat_i[22] _3715_/X _3724_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_6512_ _6510_/Y _6511_/Y _6510_/Y _6511_/Y _6545_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_147_834 VGND VPWR sky130_fd_sc_hd__decap_12
X_7492_ _7492_/HI la_data_out[19] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_174_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_558 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1118 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1227 VGND VPWR sky130_fd_sc_hd__decap_12
X_6443_ _6449_/A _6442_/X _6450_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_175_1219 VGND VPWR sky130_fd_sc_hd__fill_1
X_6374_ wbs_dat_i[2] _6364_/B _6374_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_173_196 VGND VPWR sky130_fd_sc_hd__decap_12
X_5325_ _5313_/X _5324_/X _5313_/X _5324_/X _5325_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_263 VGND VPWR sky130_fd_sc_hd__decap_12
X_5256_ _5254_/X _5255_/X _5256_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_87_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_851 VGND VPWR sky130_fd_sc_hd__decap_3
X_4207_ _4102_/Y _4104_/Y _4206_/Y _4207_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_5187_ _5178_/A _3930_/A _5187_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_112_1203 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_681 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_203 VGND VPWR sky130_fd_sc_hd__decap_8
X_4138_ _4898_/A _4137_/X _4179_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_112_1247 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_865 VGND VPWR sky130_fd_sc_hd__fill_1
X_4069_ _4038_/Y _4068_/X _4038_/Y _4068_/X _4069_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_73_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1001 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_404 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_751 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_415 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_453 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1023 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_745 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_1094 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_447 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_1059 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_648 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_727 VGND VPWR sky130_fd_sc_hd__decap_12
X_7759_ _7759_/D _5503_/A _7758_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_812 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1253 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1248 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_76 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_869 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1013 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_678 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1035 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1114 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_756 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_1158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_692 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_578 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_364 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_729 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_857 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_943 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_1142 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_879 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_1164 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_554 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_581 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_587 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_801 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_428 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_620 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_834 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_56 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_642 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_692 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_889 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_623 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_155_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1260 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1252 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1203 VGND VPWR sky130_fd_sc_hd__decap_12
X_5110_ _4547_/A _4498_/B _5110_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_174_1274 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_80 VGND VPWR sky130_fd_sc_hd__decap_12
X_6090_ _6027_/Y _6028_/B _6027_/Y _6028_/B _6090_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_33_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_147 VGND VPWR sky130_fd_sc_hd__decap_12
X_5041_ _6019_/A _6019_/B _5041_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_97_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_556 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1179 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_718 VGND VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_0_wb_clk_i wb_clk_i clkbuf_0_wb_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_20_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_898 VGND VPWR sky130_fd_sc_hd__fill_1
X_6992_ _6885_/A _6990_/Y _6991_/X _7649_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_168_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_312 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_323 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_548 VGND VPWR sky130_fd_sc_hd__fill_1
X_5943_ _5929_/X _5940_/B _5940_/X _5943_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_81_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1064 VGND VPWR sky130_fd_sc_hd__fill_2
X_5874_ _5872_/X _5873_/X _5874_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_21_401 VGND VPWR sky130_fd_sc_hd__decap_12
X_7613_ _7220_/X _7151_/A _7785_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_142_1218 VGND VPWR sky130_fd_sc_hd__decap_12
X_4825_ _4823_/X _4824_/X _4825_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_194_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_300 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_439 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_748 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1081 VGND VPWR sky130_fd_sc_hd__decap_12
X_7544_ _7544_/HI la_data_out[71] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_21_489 VGND VPWR sky130_fd_sc_hd__decap_4
X_4756_ _4589_/A _4756_/B _4756_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_175_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_333 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_653 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_269 VGND VPWR sky130_fd_sc_hd__decap_12
X_3707_ _3707_/A _3702_/X _3707_/C _3707_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_146_141 VGND VPWR sky130_fd_sc_hd__decap_12
X_4687_ _4601_/X _4602_/X _4601_/X _4602_/X _4687_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7475_ _7475_/HI la_data_out[2] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_31_1270 VGND VPWR sky130_fd_sc_hd__decap_6
X_6426_ _6421_/Y _6422_/Y _6488_/B _6426_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_179_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1038 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_550 VGND VPWR sky130_fd_sc_hd__decap_12
X_6357_ _6354_/A _6357_/B _6357_/C _6357_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_108_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_701 VGND VPWR sky130_fd_sc_hd__decap_8
X_5308_ _5128_/X _5132_/X _5131_/X _5308_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_130_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_434 VGND VPWR sky130_fd_sc_hd__decap_12
X_6288_ _5910_/X _5926_/X _5985_/A _6288_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_103_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_767 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_607 VGND VPWR sky130_fd_sc_hd__decap_12
X_5239_ _5237_/X _5238_/X _5239_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_130_575 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_151_1082 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_312 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_228 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_334 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_201 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_773 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_212 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_234 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_581 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_245 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_704 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_564 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_31 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_256 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_434 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_267 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_928 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_289 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_620 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_642 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_1094 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_450 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_664 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_984 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_770 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_420 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_347 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_829 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_572 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_165 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_850 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_489 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_1174 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1215 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1177 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_898 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1248 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_841 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_773 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_529 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_242 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1221 VGND VPWR sky130_fd_sc_hd__decap_12
X_4610_ _4608_/X _4609_/X _4813_/B VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_1005 VGND VPWR sky130_fd_sc_hd__fill_2
X_5590_ _5588_/X _5589_/X _5588_/X _5589_/X _5590_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_2090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_940 VGND VPWR sky130_fd_sc_hd__decap_12
X_4541_ _4538_/X _4539_/X _4538_/X _4539_/X _4541_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_157_973 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1049 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_983 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1189 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_239 VGND VPWR sky130_fd_sc_hd__decap_12
X_4472_ _4467_/X _4471_/X _4470_/X _4472_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_7260_ _4308_/A _7260_/B _7260_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_6211_ _6211_/A _6211_/B _6211_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_7191_ _7235_/A _7190_/X _7236_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_131_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1030 VGND VPWR sky130_fd_sc_hd__decap_12
X_6142_ _6138_/Y _6140_/X _6141_/X _7779_/D VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_112_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_851 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1085 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_776 VGND VPWR sky130_fd_sc_hd__fill_2
X_6073_ _6311_/B _6073_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_135_1066 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_426 VGND VPWR sky130_fd_sc_hd__fill_1
X_5024_ _5023_/A _5023_/B _5023_/X _5024_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_135_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_448 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_971 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6975_ _6955_/X _7019_/B _6975_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_0_1043 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_367 VGND VPWR sky130_fd_sc_hd__decap_12
X_5926_ _5911_/X _5925_/X _5926_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_62_890 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1098 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_406 VGND VPWR sky130_fd_sc_hd__decap_12
X_5857_ _5822_/X _5856_/B _5856_/Y _5857_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_179_597 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1097 VGND VPWR sky130_fd_sc_hd__fill_1
X_4808_ _4711_/X _4733_/X _4544_/X _4734_/X _4881_/A VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_210_866 VGND VPWR sky130_fd_sc_hd__decap_12
X_5788_ _3901_/X _4289_/Y _5789_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_194_556 VGND VPWR sky130_fd_sc_hd__decap_12
X_7527_ _7527_/HI la_data_out[54] VGND VPWR sky130_fd_sc_hd__conb_1
X_4739_ _4722_/X _4723_/X _4722_/X _4723_/X _4739_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_148_995 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_932 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_175_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_623 VGND VPWR sky130_fd_sc_hd__decap_12
X_7458_ _7458_/HI io_out[23] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_119_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_27 VGND VPWR sky130_fd_sc_hd__decap_12
X_6409_ _6409_/A _6409_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_134_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1130 VGND VPWR sky130_fd_sc_hd__decap_12
X_7389_ _7386_/Y _7387_/X _4812_/A _7388_/X wbs_dat_o[25] VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_116_881 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_721 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_840 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1005 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_1136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_629 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_168 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_64 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_418 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_610 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_481 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_695 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_386 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_323 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_654 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_1210 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_849 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_851 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1145 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_792 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_483 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_158_1044 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_678 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1151 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_986 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1252 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_1228 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_426 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_383 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_919 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_955 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_977 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_194 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_367 VGND VPWR sky130_fd_sc_hd__decap_12
X_6760_ _6735_/A _6735_/B _6735_/X _6759_/X _6760_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_91_1212 VGND VPWR sky130_fd_sc_hd__decap_8
X_3972_ _3952_/X _3953_/X _3952_/X _3953_/X _3972_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_204_660 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_337 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_581 VGND VPWR sky130_fd_sc_hd__decap_8
X_5711_ _5707_/X _5709_/X _5754_/A _5710_/Y _5711_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_91_1245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_6691_ _6650_/X _6689_/X _6690_/X _6691_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_149_726 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_206_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_562 VGND VPWR sky130_fd_sc_hd__decap_12
X_5642_ _5631_/X _5636_/X _5631_/X _5636_/X _5642_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_5573_ _5573_/A _5573_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_102_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1084 VGND VPWR sky130_fd_sc_hd__decap_12
X_7312_ _7312_/A _7324_/B _7312_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4524_ _4521_/X _4522_/X _4538_/B _4524_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_7243_ _7186_/X _7242_/X _6085_/X _7243_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_172_784 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_166 VGND VPWR sky130_fd_sc_hd__decap_12
X_4455_ _4455_/A _4455_/B _4456_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_160_935 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_1177 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1139 VGND VPWR sky130_fd_sc_hd__decap_12
X_4386_ _4378_/X _4382_/X _4378_/X _4382_/X _4386_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7174_ _7172_/Y _7173_/Y _7172_/Y _7173_/Y _7237_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_131_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_851 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_916 VGND VPWR sky130_fd_sc_hd__decap_12
X_6125_ _6024_/Y _6124_/X _4446_/Y _6125_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_112_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_949 VGND VPWR sky130_fd_sc_hd__decap_12
X_6056_ _6042_/A _6053_/X _6057_/C VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_85_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_779 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1252 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_1082 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_1274 VGND VPWR sky130_fd_sc_hd__decap_3
X_5007_ _4993_/X _5002_/X _4993_/X _5002_/X _5007_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_38_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_684 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1123 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_4217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_879 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_507 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_96_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_659 VGND VPWR sky130_fd_sc_hd__decap_12
X_6958_ _6956_/Y _6957_/Y _6956_/Y _6957_/Y _7021_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_3549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_849 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_39 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_11 VGND VPWR sky130_fd_sc_hd__decap_3
X_5909_ _5884_/X _5908_/X _5884_/X _5908_/X _5909_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_2848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_501 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_6889_ _6878_/X _6888_/X _6811_/X _6889_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_14_44 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_167_545 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_66 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1151 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_216 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_943 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_954 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1203 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_238 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_1225 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_784 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1119 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_968 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_309 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_702 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_724 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_41 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1038 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_1094 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_1004 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_779 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_971 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_418 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_749 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_334 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_120 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_963 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_131 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_356 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_367 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_4751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_95 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_495 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_4784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_337 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_562 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_1095 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_556 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_718 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_186_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1268 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_794 VGND VPWR sky130_fd_sc_hd__decap_12
X_4240_ _4240_/A _4240_/B _4240_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_113_147 VGND VPWR sky130_fd_sc_hd__decap_12
X_4171_ _4168_/X _4170_/X _4171_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_141_489 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_990 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_1014 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1074 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_234 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1099 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_960 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_716 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_142 VGND VPWR sky130_fd_sc_hd__decap_12
X_6812_ _6753_/X _6809_/X _6811_/X _6812_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_1_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_101 VGND VPWR sky130_fd_sc_hd__fill_1
X_7792_ _6050_/Y _7343_/A _7746_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_51_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_849 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_337 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_416 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1020 VGND VPWR sky130_fd_sc_hd__decap_12
X_6743_ la_data_in[35] _6744_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_149_501 VGND VPWR sky130_fd_sc_hd__decap_12
X_3955_ _3948_/X _3954_/X _3957_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_52_1026 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_178 VGND VPWR sky130_fd_sc_hd__decap_12
X_6674_ _6658_/X _6673_/X _6670_/X _6674_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_108_1274 VGND VPWR sky130_fd_sc_hd__decap_3
X_3886_ _5731_/A _5178_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_91_1097 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_578 VGND VPWR sky130_fd_sc_hd__fill_1
X_5625_ _4665_/A _4492_/A _5625_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_176_386 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_239 VGND VPWR sky130_fd_sc_hd__decap_12
X_5556_ _5534_/Y _5535_/X _5534_/Y _5535_/X _5556_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_191_367 VGND VPWR sky130_fd_sc_hd__decap_12
X_4507_ _4506_/A _4506_/B _4506_/X _4507_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_5487_ _4653_/A _4898_/D _5487_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_172_581 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_648 VGND VPWR sky130_fd_sc_hd__decap_12
X_7226_ _7226_/A _7194_/X _7226_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_133_968 VGND VPWR sky130_fd_sc_hd__decap_8
X_4438_ _4388_/X _4433_/X _4388_/X _4433_/X _4438_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_776 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_798 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_713 VGND VPWR sky130_fd_sc_hd__decap_12
X_7157_ _7157_/A _7157_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_116_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_510 VGND VPWR sky130_fd_sc_hd__decap_8
X_4369_ _4348_/X _4349_/X _4347_/X _4350_/X _4369_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_98_381 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_532 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_223 VGND VPWR sky130_fd_sc_hd__decap_3
X_6108_ _6095_/Y _6098_/Y _6108_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7088_ _7052_/Y _7053_/Y _7120_/B _7088_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_58_267 VGND VPWR sky130_fd_sc_hd__decap_8
X_6039_ _6038_/X _6070_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_6_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_56 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_27 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_4036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_974 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_10 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_922 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_32 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_624 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_43 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1054 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_54 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_1016 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_112 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_65 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_123 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_76 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_117 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_98 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_832 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_98 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_865 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_532 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_31 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_482 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_182_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_514 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_536 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1172 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_795 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1025 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_618 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_786 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_173_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_711 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_1151 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_206_755 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_771 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_175 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_635 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_977 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_93 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_999 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_178 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_19 _5507_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_3740_ wbs_dat_i[20] _3715_/X _3740_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_198_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_352 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_239 VGND VPWR sky130_fd_sc_hd__decap_12
X_5410_ _5200_/A _4856_/B _5410_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_173_334 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_868 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_6390_ _6390_/A _6390_/B _6390_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_127_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_902 VGND VPWR sky130_fd_sc_hd__decap_12
X_5341_ _5341_/A _4856_/B _5343_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_154_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_957 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1008 VGND VPWR sky130_fd_sc_hd__decap_12
X_5272_ _5230_/X _5251_/X _5230_/X _5251_/X _5272_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_173_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_776 VGND VPWR sky130_fd_sc_hd__decap_12
X_7011_ _6946_/X _6978_/X _7012_/C VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_87_318 VGND VPWR sky130_fd_sc_hd__decap_12
X_4223_ _4216_/X _4222_/X _4216_/X _4222_/X _4223_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_68_532 VGND VPWR sky130_fd_sc_hd__decap_12
X_4154_ _4150_/Y _4151_/X _4150_/Y _4151_/X _4200_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_210_1008 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_587 VGND VPWR sky130_fd_sc_hd__fill_1
X_4085_ _3693_/X _4126_/B _4085_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_83_524 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_790 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_1183 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1235 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_922 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1243 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_495 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_916 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_590 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_281 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_123 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_169_629 VGND VPWR sky130_fd_sc_hd__decap_12
X_7775_ _7775_/D _7775_/Q _7774_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_168_117 VGND VPWR sky130_fd_sc_hd__decap_12
X_4987_ _4986_/X _4987_/X VGND VPWR sky130_fd_sc_hd__buf_1
XPHY_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_476 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_318 VGND VPWR sky130_fd_sc_hd__decap_12
X_6726_ _6724_/Y _6725_/Y _6724_/Y _6725_/Y _6792_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_459 VGND VPWR sky130_fd_sc_hd__decap_12
X_3938_ _3938_/A _4653_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_165_813 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_852 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_824 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_684 VGND VPWR sky130_fd_sc_hd__decap_12
X_6657_ _6612_/Y _6613_/Y _6614_/X _6656_/X _6657_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_164_312 VGND VPWR sky130_fd_sc_hd__decap_12
X_3869_ _4742_/A _4718_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_137_548 VGND VPWR sky130_fd_sc_hd__fill_1
X_5608_ _5157_/A _5129_/B _5608_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_192_654 VGND VPWR sky130_fd_sc_hd__decap_12
X_6588_ _6586_/A _6539_/X _6587_/Y _6588_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_118_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_378 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_1069 VGND VPWR sky130_fd_sc_hd__decap_12
X_5539_ _5537_/X _5538_/X _5537_/X _5538_/X _5539_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_145_592 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_979 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_105_456 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_404 VGND VPWR sky130_fd_sc_hd__fill_1
X_7209_ _7144_/X _7203_/B _7209_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_191_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_489 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_543 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1059 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_220 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_635 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_202 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_977 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_145 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_426 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_769 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_638 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_971 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1182 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_852 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_801 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_846 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_323 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_334 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_548 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_155_356 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_367 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_196_1158 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_529 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_581 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_540 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_562 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_595 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_437 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_971 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_1085 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_395 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_708 VGND VPWR sky130_fd_sc_hd__decap_12
X_4910_ _4900_/X _4909_/X _4900_/X _4909_/X _4910_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_92_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_549 VGND VPWR sky130_fd_sc_hd__decap_4
X_5890_ _5887_/X _5888_/X _5889_/X _5890_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_209_1224 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_916 VGND VPWR sky130_fd_sc_hd__decap_12
X_4841_ _4841_/A _4915_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_179_949 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_774 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_999 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_178_459 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_1170 VGND VPWR sky130_fd_sc_hd__decap_12
X_7560_ _7560_/HI la_data_out[87] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_53_1132 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1252 VGND VPWR sky130_fd_sc_hd__decap_12
X_4772_ _4772_/A _4771_/X _4772_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_147_802 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_1105 VGND VPWR sky130_fd_sc_hd__decap_12
X_6511_ la_data_in[8] _6511_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_3723_ _4539_/A _3712_/X _3725_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_159_684 VGND VPWR sky130_fd_sc_hd__decap_12
X_7491_ _7491_/HI la_data_out[18] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_174_621 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_526 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_846 VGND VPWR sky130_fd_sc_hd__decap_8
X_6442_ _6387_/A _6387_/B _6387_/X _6441_/X _6442_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_174_654 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_162_816 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_134_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_161_315 VGND VPWR sky130_fd_sc_hd__decap_8
X_6373_ _4898_/D _6373_/B _6375_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_161_326 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_0_0_wb_clk_i clkbuf_2_0_1_wb_clk_i/X clkbuf_3_0_0_wb_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_5324_ _5322_/X _5323_/X _5322_/X _5323_/X _5324_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_88_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_916 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_509 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_938 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_798 VGND VPWR sky130_fd_sc_hd__fill_1
X_5255_ _4665_/A _4299_/X _5255_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4206_ _4206_/A _4206_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_102_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_863 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_1234 VGND VPWR sky130_fd_sc_hd__decap_12
X_5186_ _5186_/A _4743_/B _5186_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_96_660 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_971 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_362 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_1136 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_373 VGND VPWR sky130_fd_sc_hd__decap_12
X_4137_ _4460_/B _4137_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_96_693 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_215 VGND VPWR sky130_fd_sc_hd__fill_2
X_4068_ _4065_/X _4067_/B _4067_/X _4068_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_3_1052 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_933 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_405 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_416 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_977 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_426 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_1035 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_757 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_273 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_459 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_1221 VGND VPWR sky130_fd_sc_hd__decap_4
X_7758_ _7758_/D _5632_/A _7758_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_739 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6709_ _6709_/A _6709_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_119 VGND VPWR sky130_fd_sc_hd__decap_3
X_7689_ _7689_/D _7689_/Q _7707_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_22_44 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_193_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_837 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1150 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1172 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_156_1142 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1126 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_971 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_513 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_524 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_481 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_877 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_376 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1176 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_62 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_1135 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_1266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_413 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_245 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_593 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_813 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_457 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_312 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_660 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_632 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_846 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_68 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_654 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_849 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1130 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1212 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1272 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_679 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1215 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_1158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_881 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_1237 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_392 VGND VPWR sky130_fd_sc_hd__decap_12
X_5040_ _5040_/A _6019_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_111_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_568 VGND VPWR sky130_fd_sc_hd__decap_12
X_6991_ la_data_in[79] _6991_/B _6991_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_0_1203 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_1142 VGND VPWR sky130_fd_sc_hd__decap_12
X_5942_ _5911_/X _5925_/X _5926_/X _5942_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_80_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_240 VGND VPWR sky130_fd_sc_hd__decap_4
X_5873_ _5830_/X _5837_/X _5830_/X _5837_/X _5873_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_34_785 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1246 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_413 VGND VPWR sky130_fd_sc_hd__decap_12
X_7612_ _7612_/D _7154_/A _7729_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_22_947 VGND VPWR sky130_fd_sc_hd__decap_12
X_4824_ _4824_/A _4492_/A _4824_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_166_407 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_727 VGND VPWR sky130_fd_sc_hd__decap_8
X_7543_ _7543_/HI la_data_out[70] VGND VPWR sky130_fd_sc_hd__conb_1
X_4755_ _4631_/B _4756_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_18_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_952 VGND VPWR sky130_fd_sc_hd__decap_12
X_3706_ wbs_adr_i[30] _3706_/B _3704_/X _3705_/X _3707_/C VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_119_345 VGND VPWR sky130_fd_sc_hd__decap_12
X_7474_ _7474_/HI la_data_out[1] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_147_665 VGND VPWR sky130_fd_sc_hd__decap_6
X_4686_ _4677_/X _4683_/X _4684_/X _4685_/X _4686_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_179_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_827 VGND VPWR sky130_fd_sc_hd__fill_1
X_6425_ _6487_/A _6487_/B _6488_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_49_1009 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_123 VGND VPWR sky130_fd_sc_hd__decap_12
X_6356_ wbs_dat_i[7] _6349_/B _6357_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_115_562 VGND VPWR sky130_fd_sc_hd__decap_12
X_5307_ _4769_/X _4773_/X _4769_/X _4773_/X _5307_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_103_724 VGND VPWR sky130_fd_sc_hd__decap_8
X_6287_ _6219_/X _6285_/X _6286_/X _6287_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_130_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_757 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_446 VGND VPWR sky130_fd_sc_hd__decap_12
X_5238_ _5215_/X _5216_/X _5217_/X _5238_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_103_779 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_619 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_660 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_68 VGND VPWR sky130_fd_sc_hd__decap_12
X_5169_ _4678_/A _4747_/B _5169_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_111_790 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_630 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_151_1094 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_708 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1067 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_1007 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_346 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_140_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_99 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_202 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_903 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_213 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_785 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_224 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_158_919 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_593 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_257 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_268 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_576 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_446 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_279 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_417 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1024 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_149_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_490 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_462 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_782 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_624 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_432 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_668 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_359 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_165_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_177 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_595 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_862 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_603 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1186 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_663 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1189 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_590 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_853 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_785 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_582 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_886 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_727 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_254 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_952 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_1203 VGND VPWR sky130_fd_sc_hd__decap_12
X_4540_ _4540_/A _4540_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1157 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_922 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_35 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_995 VGND VPWR sky130_fd_sc_hd__decap_12
X_4471_ _4470_/A _4469_/X _4470_/X _4471_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_183_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_337 VGND VPWR sky130_fd_sc_hd__decap_12
X_6210_ _6219_/A _6202_/B _6209_/Y _4540_/A _6109_/X _6211_/B VGND VPWR sky130_fd_sc_hd__a32oi_4
XFILLER_116_359 VGND VPWR sky130_fd_sc_hd__decap_12
X_7190_ _7172_/Y _7173_/Y _7238_/B _7190_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_48_1020 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_318 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_1042 VGND VPWR sky130_fd_sc_hd__decap_6
X_6141_ _4248_/Y _6103_/X _6092_/X _6141_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_112_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_755 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1097 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_863 VGND VPWR sky130_fd_sc_hd__decap_12
X_6072_ _3967_/X _6072_/B _6072_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_57_107 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1078 VGND VPWR sky130_fd_sc_hd__decap_12
X_5023_ _5023_/A _5023_/B _5023_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_39_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_983 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1022 VGND VPWR sky130_fd_sc_hd__fill_1
X_6974_ _6956_/Y _6957_/Y _7022_/B _7019_/B VGND VPWR sky130_fd_sc_hd__o21a_4
XPHY_3709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_1191 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_1040 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1160 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1055 VGND VPWR sky130_fd_sc_hd__decap_12
X_5925_ _5912_/X _5922_/X _5923_/X _5924_/X _5925_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_80_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_593 VGND VPWR sky130_fd_sc_hd__fill_1
X_5856_ _5822_/X _5856_/B _5856_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_16_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_716 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_418 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_1136 VGND VPWR sky130_fd_sc_hd__decap_12
X_4807_ _4806_/A _4806_/B _4806_/Y _4807_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_166_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_788 VGND VPWR sky130_fd_sc_hd__decap_4
X_5787_ _5787_/A _4901_/A _5789_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_210_878 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_194_568 VGND VPWR sky130_fd_sc_hd__decap_12
X_7526_ _7526_/HI la_data_out[53] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_147_440 VGND VPWR sky130_fd_sc_hd__decap_12
X_4738_ _4725_/X _4726_/X _4725_/X _4726_/X _4738_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_163_900 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_410 VGND VPWR sky130_fd_sc_hd__decap_12
X_7457_ _7457_/HI io_out[22] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_135_635 VGND VPWR sky130_fd_sc_hd__decap_12
X_4669_ _4666_/X _4667_/X _4668_/X _4669_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_163_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_6408_ _6408_/A _6408_/B _6408_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_123_819 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_605 VGND VPWR sky130_fd_sc_hd__decap_8
X_7388_ _7388_/A _7388_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_134_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_638 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_626 VGND VPWR sky130_fd_sc_hd__decap_8
X_6339_ _6350_/A _6337_/X _6339_/C _6339_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_118_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_637 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_648 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_153_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_125 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_852 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_863 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_140 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_76 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_471 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_622 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_493 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_398 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_357 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_508 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_1222 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_863 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_530 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_727 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1119 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_513 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_788 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_265 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_546 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_197_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_954 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_999 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_1163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_153_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1174 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1231 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_998 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1212 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_841 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_874 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_395 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_967 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_184 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_806 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_1038 VGND VPWR sky130_fd_sc_hd__decap_12
X_3971_ _3948_/X _3954_/X _3970_/Y _3971_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_5710_ _5707_/X _5709_/X _5707_/X _5709_/X _5710_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_50_349 VGND VPWR sky130_fd_sc_hd__decap_12
X_6690_ _6670_/A _6690_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_93_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_885 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_5641_ _5637_/X _5638_/X _5639_/Y _5640_/X _5641_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_31_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_557 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_440 VGND VPWR sky130_fd_sc_hd__decap_12
X_5572_ _5561_/X _5562_/X _5561_/X _5562_/X _5572_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_106_1180 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_1191 VGND VPWR sky130_fd_sc_hd__decap_8
X_7311_ io_in[14] _7312_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_4523_ _4521_/X _4522_/X _4538_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_144_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1044 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1096 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_145_977 VGND VPWR sky130_fd_sc_hd__decap_12
X_7242_ _7604_/Q la_data_in[98] _7180_/X _7242_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_105_819 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1028 VGND VPWR sky130_fd_sc_hd__decap_8
X_4454_ _4655_/A _4748_/B _4456_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_132_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_796 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_1189 VGND VPWR sky130_fd_sc_hd__fill_1
X_7173_ la_data_in[100] _7173_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4385_ _4322_/Y _4384_/Y _4385_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_131_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_552 VGND VPWR sky130_fd_sc_hd__decap_12
X_6124_ _4450_/X _4451_/X _6124_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_86_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_928 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_671 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_373 VGND VPWR sky130_fd_sc_hd__decap_12
X_6055_ _7338_/A _6059_/B _6055_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_105_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_546 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_257 VGND VPWR sky130_fd_sc_hd__decap_12
X_5006_ _5003_/Y _5005_/B _5005_/X _5006_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_82_920 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_471 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1067 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_110 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_335 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_452 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6957_ la_data_in[68] _6957_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_3539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5908_ _5885_/X _5905_/X _5906_/X _5907_/X _5908_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XPHY_2838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6888_ _6822_/A la_data_in[61] _6824_/X _6888_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XPHY_2849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_703 VGND VPWR sky130_fd_sc_hd__decap_12
X_5839_ _5825_/X _5839_/B _5839_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_14_78 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_708 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_771 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_398 VGND VPWR sky130_fd_sc_hd__decap_12
X_7509_ _7509_/HI la_data_out[36] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_175_590 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_646 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_966 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_120_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_44 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1237 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_714 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_53 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_728 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_162 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_825 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_1167 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_403 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_806 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_206_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_143 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_154 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_305 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_189_159 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_658 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1052 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1022 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_199_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1066 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1099 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_782 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1258 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_468 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_703 VGND VPWR sky130_fd_sc_hd__decap_4
X_4170_ _4919_/A _4591_/B _4170_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_110_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_171_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_972 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_728 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_419 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_471 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_633 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_208_285 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_666 VGND VPWR sky130_fd_sc_hd__decap_12
X_6811_ _6905_/A _6811_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_91_772 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_154 VGND VPWR sky130_fd_sc_hd__decap_12
X_7791_ _6057_/X _7338_/A _7785_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_1_1172 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_794 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_196_608 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_647 VGND VPWR sky130_fd_sc_hd__decap_12
X_6742_ _6742_/A _6744_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_3954_ _3952_/X _3953_/X _3951_/X _3954_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_211_428 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_1032 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_1111 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_1163 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_861 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1171 VGND VPWR sky130_fd_sc_hd__decap_12
X_6673_ _7694_/Q la_data_in[28] _6608_/X _6673_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_3885_ _7796_/Q _5731_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_17_1158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_708 VGND VPWR sky130_fd_sc_hd__decap_8
X_5624_ _5623_/A _5622_/X _5623_/X _5624_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_164_505 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_1128 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_858 VGND VPWR sky130_fd_sc_hd__decap_12
X_5555_ _5310_/X _5311_/X _5299_/X _5312_/X _5555_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_145_730 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_903 VGND VPWR sky130_fd_sc_hd__decap_12
X_4506_ _4506_/A _4506_/B _4506_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_191_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_251 VGND VPWR sky130_fd_sc_hd__decap_12
X_5486_ _4548_/A _4778_/B _5486_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_160_711 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_936 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_487 VGND VPWR sky130_fd_sc_hd__fill_1
X_7225_ _7210_/A _7225_/B _7224_/Y _7225_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_4437_ _4434_/Y _4436_/B _4436_/X _4437_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_28_1210 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1123 VGND VPWR sky130_fd_sc_hd__decap_12
X_7156_ _7154_/Y _7155_/Y _7156_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_132_479 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_660 VGND VPWR sky130_fd_sc_hd__decap_8
X_4368_ _4368_/A _4368_/B _4368_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_59_725 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_202 VGND VPWR sky130_fd_sc_hd__decap_12
X_6107_ _6095_/A _6097_/X _6107_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_98_393 VGND VPWR sky130_fd_sc_hd__decap_4
X_7087_ _7119_/A _7119_/B _7120_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_101_855 VGND VPWR sky130_fd_sc_hd__decap_12
X_4299_ _4569_/B _4299_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_86_555 VGND VPWR sky130_fd_sc_hd__decap_12
X_6038_ _6038_/A _6038_/B wbs_we_i _7261_/A _6038_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_27_611 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_622 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_132_68 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_441 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1011 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_11 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_997 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_154 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_33 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_44 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_934 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_636 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_55 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1066 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_66 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1028 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_293 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_77 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_135 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_88 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_129 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_844 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_962 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_371 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_877 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_900 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_899 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_43 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_494 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_869 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_548 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_508 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1067 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_766 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_798 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_503 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_536 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_227 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_2_0_wb_clk_i clkbuf_4_3_0_wb_clk_i/A _7624_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_73_783 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_688 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_794 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_422 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_162_1008 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_647 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_861 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_158_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_346 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1044 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_763 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_1172 VGND VPWR sky130_fd_sc_hd__decap_12
X_5340_ _5185_/A _4852_/B _5340_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_115_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_142_711 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_154_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_284 VGND VPWR sky130_fd_sc_hd__decap_3
X_5271_ _5267_/X _5270_/X _5267_/X _5270_/X _5271_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_115_969 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_446 VGND VPWR sky130_fd_sc_hd__decap_12
X_7010_ _6913_/A _7012_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_4222_ _4220_/X _4221_/X _4219_/X _4222_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_142_788 VGND VPWR sky130_fd_sc_hd__decap_12
X_4153_ _4109_/X _4152_/X _4153_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_110_630 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_853 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_886 VGND VPWR sky130_fd_sc_hd__decap_12
X_4084_ _4081_/X _4082_/X _4083_/X _4086_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_55_216 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_536 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1203 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_1195 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_761 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1274 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_934 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_411 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_619 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_939 VGND VPWR sky130_fd_sc_hd__decap_12
X_4986_ _4986_/A _4985_/X _4986_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7774_ _6173_/Y _7774_/Q _7774_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_129 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3937_ _4664_/A _3938_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_6725_ la_data_in[41] _6725_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_149_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1083 VGND VPWR sky130_fd_sc_hd__decap_12
X_6656_ _6615_/Y _6616_/Y _6655_/X _6656_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_3868_ _3867_/Y _4742_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_165_836 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_886 VGND VPWR sky130_fd_sc_hd__decap_12
X_5607_ _5348_/A _4903_/B _5607_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_191_110 VGND VPWR sky130_fd_sc_hd__decap_12
X_6587_ _6524_/X _6539_/B _6587_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_3799_ _3759_/A _3822_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_192_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_903 VGND VPWR sky130_fd_sc_hd__decap_12
X_5538_ _4794_/Y _4795_/X _4794_/Y _4795_/X _5538_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1218 VGND VPWR sky130_fd_sc_hd__fill_2
X_5469_ _5467_/X _5468_/X _5469_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_87_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_7208_ _7404_/A _7206_/Y _7207_/X _7617_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_132_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_831 VGND VPWR sky130_fd_sc_hd__decap_12
X_7139_ _7210_/A _7139_/B _7138_/Y _7139_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_154_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_330 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_555 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_189_1111 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_566 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1005 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_1189 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_189_1144 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_290 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_463 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_160_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_76 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_794 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_647 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_764 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1000 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1041 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_983 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_825 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_864 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_813 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_858 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_184 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_806 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_182_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_711 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_349 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_606 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_540 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_551 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_449 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_801 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1097 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1228 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_206_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_506 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_761 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_1203 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_528 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_956 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_928 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_1236 VGND VPWR sky130_fd_sc_hd__decap_3
X_4840_ _4639_/X _4643_/X _4642_/X _4840_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XPHY_4390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_786 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1111 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_477 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_4771_ _4771_/A _4570_/B _4771_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_194_909 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_1182 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_1144 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1264 VGND VPWR sky130_fd_sc_hd__decap_12
X_6510_ _6510_/A _6510_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_3722_ _3722_/A _4539_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_7490_ _7490_/HI la_data_out[17] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_14_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_633 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_538 VGND VPWR sky130_fd_sc_hd__decap_8
X_6441_ _6390_/A _6390_/B _6390_/X _6440_/X _6441_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_140_1158 VGND VPWR sky130_fd_sc_hd__decap_12
X_6372_ _6381_/A _6372_/B _6371_/Y _7733_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_161_338 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_733 VGND VPWR sky130_fd_sc_hd__decap_8
X_5323_ _5183_/X _5193_/X _5168_/X _5194_/X _5323_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_115_755 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_617 VGND VPWR sky130_fd_sc_hd__decap_12
X_5254_ _4678_/A _4293_/X _5254_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_114_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_831 VGND VPWR sky130_fd_sc_hd__decap_12
X_4205_ _4211_/B _4205_/B _6027_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_151_1221 VGND VPWR sky130_fd_sc_hd__decap_12
X_5185_ _5185_/A _3938_/A _5185_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_25_1246 VGND VPWR sky130_fd_sc_hd__decap_4
X_4136_ _4757_/B _4460_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_110_471 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_547 VGND VPWR sky130_fd_sc_hd__fill_1
X_4067_ _4065_/X _4067_/B _4067_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_3_1042 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1064 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_1071 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1097 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_1044 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_945 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_406 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_417 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_196_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_764 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_769 VGND VPWR sky130_fd_sc_hd__decap_12
X_4969_ _4929_/X _4930_/X _4928_/X _4931_/X _4969_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_7757_ _7757_/D _5639_/A _7756_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6708_ _6694_/X _6705_/A _6707_/X _7682_/D VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_138_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_23 VGND VPWR sky130_fd_sc_hd__decap_8
X_7688_ _6692_/X _6624_/A _7707_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_32_1228 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_324 VGND VPWR sky130_fd_sc_hd__fill_1
X_6639_ _7683_/Q _6639_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_192_441 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_964 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_593 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_1121 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_541 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1138 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_650 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_20 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_983 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_807 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_536 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_867 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_889 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_772 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_388 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_783 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_455 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_1245 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1008 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_1188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_263 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_425 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_959 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_471 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_129_825 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_791 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_672 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_666 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_368 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_891 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1224 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_937 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_596 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1249 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_257 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1148 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_141 VGND VPWR sky130_fd_sc_hd__decap_12
X_6990_ la_data_in[79] _6991_/B _6990_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_25_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_697 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_1154 VGND VPWR sky130_fd_sc_hd__decap_12
X_5941_ _5928_/X _5940_/X _5928_/X _5938_/X _5941_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_19_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_361 VGND VPWR sky130_fd_sc_hd__decap_12
X_5872_ _5870_/X _5871_/X _5872_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_178_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_764 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_550 VGND VPWR sky130_fd_sc_hd__decap_12
X_4823_ _4822_/A _4821_/X _4887_/A _4823_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_7611_ _7225_/X _7157_/A _7729_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_21_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_1099 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_458 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1061 VGND VPWR sky130_fd_sc_hd__decap_6
X_4754_ _4740_/X _4746_/X _4752_/X _4753_/X _4754_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_7542_ _7542_/HI la_data_out[69] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_147_611 VGND VPWR sky130_fd_sc_hd__fill_2
X_3705_ wbs_adr_i[20] wbs_adr_i[23] wbs_adr_i[22] wbs_adr_i[25] _3705_/X VGND VPWR
+ sky130_fd_sc_hd__or4_4
X_7473_ _7473_/HI la_data_out[0] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_175_964 VGND VPWR sky130_fd_sc_hd__decap_12
X_4685_ _4677_/X _4683_/X _4677_/X _4683_/X _4685_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_119_357 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1154 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_119_379 VGND VPWR sky130_fd_sc_hd__decap_4
X_6424_ _6421_/Y _6422_/Y _6421_/Y _6422_/Y _6487_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_108_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_349 VGND VPWR sky130_fd_sc_hd__decap_12
X_6355_ _4346_/B _6348_/B _6357_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_89_904 VGND VPWR sky130_fd_sc_hd__decap_8
X_5306_ _5303_/X _5304_/X _5532_/B _5306_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_143_883 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_574 VGND VPWR sky130_fd_sc_hd__decap_12
X_6286_ _5807_/Y _6216_/X _3743_/A _6286_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_102_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_329 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_544 VGND VPWR sky130_fd_sc_hd__decap_12
X_5237_ _5232_/X _5236_/X _5232_/X _5236_/X _5237_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_9_1262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1032 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_588 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1054 VGND VPWR sky130_fd_sc_hd__decap_8
X_5168_ _5154_/X _5167_/X _5154_/X _5167_/X _5168_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_151_1062 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_525 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_1024 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_642 VGND VPWR sky130_fd_sc_hd__decap_12
X_4119_ _5304_/A _4164_/B _4119_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_5099_ _5099_/A _4906_/B _5099_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_204_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1019 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_528 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_83_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_753 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_68 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_203 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_701 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_225 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_263 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_236 VGND VPWR sky130_fd_sc_hd__decap_3
X_7809_ _3783_/Y _7809_/Q _7806_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_247 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_257 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_269 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_588 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_600 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1052 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_789 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_429 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_162_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_99 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_603 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_1205 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_474 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_636 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1249 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_444 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_872 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_393 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_615 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_791 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_631 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_845 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1198 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_601 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_506 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_1228 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_810 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_678 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_865 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_611 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_622 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_266 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1245 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_288 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_761 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_440 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1169 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_997 VGND VPWR sky130_fd_sc_hd__decap_12
X_4470_ _4470_/A _4469_/X _4470_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_117_839 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_422 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_183_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_349 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_144_669 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_701 VGND VPWR sky130_fd_sc_hd__fill_1
X_6140_ _6138_/A _6137_/X _6319_/C _6140_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_139_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_544 VGND VPWR sky130_fd_sc_hd__decap_8
X_6071_ _6317_/C _6256_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_140_875 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_717 VGND VPWR sky130_fd_sc_hd__decap_12
X_5022_ _5020_/Y _5021_/X _5020_/Y _5021_/X _5023_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_85_428 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_491 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_506 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_995 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1001 VGND VPWR sky130_fd_sc_hd__fill_2
X_6973_ _7021_/A _7021_/B _7022_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_65_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1090 VGND VPWR sky130_fd_sc_hd__decap_8
X_5924_ _5912_/X _5922_/X _5912_/X _5922_/X _5924_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_1052 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1067 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_179_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_1036 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_802 VGND VPWR sky130_fd_sc_hd__decap_12
X_5855_ _5823_/X _5852_/X _5853_/X _5854_/X _5856_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_142_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_391 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_167_728 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_181_1077 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_1148 VGND VPWR sky130_fd_sc_hd__decap_8
X_4806_ _4806_/A _4806_/B _4806_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_166_227 VGND VPWR sky130_fd_sc_hd__decap_12
X_5786_ _5178_/A _4363_/A _5786_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_119_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_277 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_15_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/X _7774_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_7525_ _7525_/HI la_data_out[52] VGND VPWR sky130_fd_sc_hd__conb_1
X_4737_ _4728_/X _4729_/X _4728_/X _4729_/X _4737_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_147_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_912 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_794 VGND VPWR sky130_fd_sc_hd__decap_12
X_4668_ _4666_/X _4667_/X _4668_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7456_ _7456_/HI io_out[21] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_162_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_647 VGND VPWR sky130_fd_sc_hd__decap_12
X_6407_ la_data_in[118] _6408_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_190_764 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1110 VGND VPWR sky130_fd_sc_hd__decap_12
X_4599_ _4596_/X _4597_/X _4598_/X _4599_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_7387_ _7387_/A _7387_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_6338_ wbs_dat_i[12] _6338_/B _6339_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_66_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_137 VGND VPWR sky130_fd_sc_hd__fill_2
X_6269_ _6269_/A _6269_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_95_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_44 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_88 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_634 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1250 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1234 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1204 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_520 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_875 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_745 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_198_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_542 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_739 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_255 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_20 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_558 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_201_1103 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_139_997 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1062 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_809 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_850 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_966 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_180_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_628 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1186 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1243 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1265 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_853 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1249 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_886 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_428 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_693 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1120 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_623 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_837 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_1036 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_859 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_169_1197 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_818 VGND VPWR sky130_fd_sc_hd__decap_12
X_3970_ _3957_/A _3970_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_62_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_486 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_897 VGND VPWR sky130_fd_sc_hd__decap_12
X_5640_ _5637_/X _5638_/X _5637_/X _5638_/X _5640_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_188_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_586 VGND VPWR sky130_fd_sc_hd__decap_12
X_5571_ _5567_/X _5568_/X _5569_/X _5570_/X _5573_/A VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_176_569 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_208 VGND VPWR sky130_fd_sc_hd__decap_12
X_4522_ _3738_/A _4565_/B _4522_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7310_ _7310_/A _7292_/B _7310_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_8_771 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_144_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_281 VGND VPWR sky130_fd_sc_hd__decap_12
X_4453_ _4453_/A _4655_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_7241_ _7187_/X _7239_/X _7240_/Y _7241_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_172_764 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_308 VGND VPWR sky130_fd_sc_hd__fill_1
X_7172_ _7606_/Q _7172_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4384_ _4383_/X _4384_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_98_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_691 VGND VPWR sky130_fd_sc_hd__decap_4
X_6123_ _4317_/X _6123_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_124_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_564 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_683 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_27 VGND VPWR sky130_fd_sc_hd__decap_12
X_6054_ _6053_/X _6059_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_140_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1221 VGND VPWR sky130_fd_sc_hd__decap_12
X_5005_ _5003_/Y _5005_/B _5005_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_100_558 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_781 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_94_792 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_932 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_121_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_105 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1248 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_464 VGND VPWR sky130_fd_sc_hd__decap_12
X_6956_ _7638_/Q _6956_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_121_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_306 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_330 VGND VPWR sky130_fd_sc_hd__decap_12
X_5907_ _5901_/X _5902_/X _5896_/X _5903_/X _5907_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XPHY_2828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_520 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6887_ _6912_/A _6880_/X _6886_/Y _6887_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_194_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_385 VGND VPWR sky130_fd_sc_hd__fill_1
X_5838_ _5826_/X _5829_/X _5830_/X _5837_/X _5839_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_10_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_895 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_889 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_1191 VGND VPWR sky130_fd_sc_hd__decap_8
X_5769_ _5655_/X _5662_/X _5654_/X _5663_/X _5769_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_148_783 VGND VPWR sky130_fd_sc_hd__decap_12
X_7508_ _7508_/HI la_data_out[35] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_108_625 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_1178 VGND VPWR sky130_fd_sc_hd__decap_12
X_7439_ io_oeb[34] _7439_/LO VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_190_550 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_606 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_1249 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_162_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_572 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_200_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_937 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_958 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_118_1030 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_672 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_417 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_461 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_415 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_818 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_44_166 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_317 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_531 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_812 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1034 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_1045 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1078 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_1215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_444 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_306 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_403 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1013 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_834 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_601 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_765 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_483 VGND VPWR sky130_fd_sc_hd__decap_12
X_6810_ wb_rst_i _6905_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_208_297 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_678 VGND VPWR sky130_fd_sc_hd__decap_12
X_7790_ _6059_/Y _7332_/A _7746_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_91_784 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1184 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_1180 VGND VPWR sky130_fd_sc_hd__decap_8
X_6741_ _6739_/Y _6740_/Y _6739_/Y _6740_/Y _6741_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_3953_ _4535_/A _4164_/B _3953_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_56_1142 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_993 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_391 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_176_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1175 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1183 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_873 VGND VPWR sky130_fd_sc_hd__decap_12
X_3884_ _3866_/X _3884_/B _3884_/C _7797_/D VGND VPWR sky130_fd_sc_hd__nor3_4
X_6672_ _6659_/X _6669_/X _6671_/Y _6672_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_143_1167 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1099 VGND VPWR sky130_fd_sc_hd__decap_12
X_5623_ _5623_/A _5622_/X _5623_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_164_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_837 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_923 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_934 VGND VPWR sky130_fd_sc_hd__decap_12
X_5554_ _5293_/X _5294_/X _5292_/Y _5295_/X _5554_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_145_742 VGND VPWR sky130_fd_sc_hd__decap_12
X_4505_ _4505_/A _4505_/B _4506_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_5485_ _5480_/X _5484_/X _5483_/X _5485_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_144_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_80 VGND VPWR sky130_fd_sc_hd__decap_12
X_4436_ _4434_/Y _4436_/B _4436_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7224_ _7224_/A _7224_/B _7224_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_116_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1222 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_609 VGND VPWR sky130_fd_sc_hd__fill_1
X_4367_ _4360_/X _4366_/X _4359_/X _4368_/B VGND VPWR sky130_fd_sc_hd__o21a_4
X_7155_ la_data_in[106] _7155_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_154_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_1135 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1266 VGND VPWR sky130_fd_sc_hd__decap_8
X_6106_ _6311_/B _6106_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_63_1168 VGND VPWR sky130_fd_sc_hd__fill_1
X_7086_ _7057_/A _7057_/B _7057_/X _7085_/X _7119_/B VGND VPWR sky130_fd_sc_hd__o22a_4
X_4298_ _4613_/B _4569_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_115_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_867 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_86_567 VGND VPWR sky130_fd_sc_hd__decap_12
X_6037_ _3710_/A _7264_/A _7261_/A VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_4005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_403 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_1023 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_453 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_3304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_604 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_23 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_166 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_34 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_67 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6939_ la_data_in[74] _6940_/B VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_3359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_78 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_89 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_812 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_147 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_171 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_856 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_1128 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_211_974 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_383 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_462 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_194_141 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_127_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_686 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_912 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_55 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_202_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_383 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_236 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_515 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_1090 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_111 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_291 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_924 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_205_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_80 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_609 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_659 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_300 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_873 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_963 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_186_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_517 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_173_314 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_528 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_775 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1146 VGND VPWR sky130_fd_sc_hd__decap_12
X_5270_ _5268_/X _5269_/X _5268_/X _5269_/X _5270_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_181_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_147 VGND VPWR sky130_fd_sc_hd__decap_12
X_4221_ _3773_/X _4328_/B _4221_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4152_ _4110_/X _4149_/X _4150_/Y _4151_/X _4152_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_110_642 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_865 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_556 VGND VPWR sky130_fd_sc_hd__decap_12
X_4083_ _4081_/X _4082_/X _4083_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_96_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_943 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_1166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_784 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_609 VGND VPWR sky130_fd_sc_hd__fill_1
X_7773_ _7773_/D _7773_/Q _7774_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4985_ _4877_/X _4878_/X _4809_/X _4879_/X _4985_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XPHY_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6724_ _7675_/Q _6724_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_189_480 VGND VPWR sky130_fd_sc_hd__decap_8
X_3936_ _7743_/Q _4664_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_108_1051 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_681 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_141 VGND VPWR sky130_fd_sc_hd__decap_12
X_6655_ _6617_/X _6654_/X _6655_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_3867_ _3867_/A _3867_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_109_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1095 VGND VPWR sky130_fd_sc_hd__decap_12
X_5606_ _5137_/A _4906_/B _5606_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_165_848 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_898 VGND VPWR sky130_fd_sc_hd__decap_12
X_6586_ _6586_/A _6541_/X _6585_/Y _6586_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_3798_ _4467_/A _3798_/B _3798_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_192_678 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_550 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_764 VGND VPWR sky130_fd_sc_hd__decap_12
X_5537_ _5526_/X _5527_/X _5525_/X _5528_/X _5537_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_106_915 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_926 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_712 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_160_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_959 VGND VPWR sky130_fd_sc_hd__decap_12
X_5468_ _5234_/A _4915_/B _5468_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7207_ la_data_in[111] _7207_/B _7207_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_4419_ _4368_/A _4368_/B _4368_/X _4419_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_99_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_501 VGND VPWR sky130_fd_sc_hd__decap_12
X_5399_ _5389_/X _5390_/X _5389_/X _5390_/X _5399_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_692 VGND VPWR sky130_fd_sc_hd__decap_12
X_7138_ _7077_/A _7138_/B _7138_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_101_620 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_843 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_631 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_578 VGND VPWR sky130_fd_sc_hd__decap_12
X_7069_ _7067_/Y _7068_/Y _7069_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_115_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1156 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_44 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_475 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_710 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_88 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_3134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_153_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_659 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_215 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_428 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_467 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1012 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_489 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_32 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1053 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_331 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_995 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_876 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_825 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_313 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_1138 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_723 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_163_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1010 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_574 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_428 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_854 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_813 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_526 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_932 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_868 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_968 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_607 VGND VPWR sky130_fd_sc_hd__decap_3
X_4770_ _4514_/A _4569_/B _4772_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_159_631 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_798 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_489 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_117 VGND VPWR sky130_fd_sc_hd__decap_12
X_3721_ _4565_/A _3722_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_158_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1156 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_151 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_483 VGND VPWR sky130_fd_sc_hd__decap_3
X_6440_ _6391_/Y _6393_/B _6393_/X _6439_/X _6440_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_127_550 VGND VPWR sky130_fd_sc_hd__decap_12
X_6371_ wbs_dat_i[3] _6364_/B _6371_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_5322_ _5318_/X _5321_/X _5318_/X _5321_/X _5322_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_142_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1093 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_767 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_907 VGND VPWR sky130_fd_sc_hd__decap_8
X_5253_ _5602_/A _4366_/B _5253_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_130_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_821 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_1200 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1252 VGND VPWR sky130_fd_sc_hd__decap_12
X_4204_ _4153_/X _4202_/X _4203_/X _4205_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_138_1099 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_843 VGND VPWR sky130_fd_sc_hd__decap_8
X_5184_ _5176_/X _5180_/X _5176_/X _5180_/X _5184_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_151_1233 VGND VPWR sky130_fd_sc_hd__decap_4
X_4135_ _4277_/A _4757_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_84_835 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_27 VGND VPWR sky130_fd_sc_hd__decap_12
X_4066_ _3998_/X _4025_/X _4026_/X _4067_/B VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_83_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_1050 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_184_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1083 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_957 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_220 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_407 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_418 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_428 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1201 VGND VPWR sky130_fd_sc_hd__decap_12
X_7756_ _7756_/D _5754_/A _7756_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4968_ _4403_/X _4404_/X _4403_/X _4404_/X _4968_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6707_ _6641_/A la_data_in[16] _6707_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1245 VGND VPWR sky130_fd_sc_hd__decap_8
X_3919_ _3919_/A _4648_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_178_984 VGND VPWR sky130_fd_sc_hd__fill_1
X_7687_ _6696_/X _6627_/A _7658_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4899_ _4949_/B _4900_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_138_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_623 VGND VPWR sky130_fd_sc_hd__decap_12
X_6638_ _6636_/Y _6638_/B _6638_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_149_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_453 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_68 VGND VPWR sky130_fd_sc_hd__decap_12
X_6569_ _6549_/X _6568_/X _6481_/X _6569_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_118_572 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_662 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_684 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_819 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_995 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_849 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_795 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_261 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_916 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_748 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_927 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_489 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_437 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_269 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_459 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_910 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_590 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_611 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_150 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_453 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_154 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1116 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1236 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_850 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_861 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_504 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_367 VGND VPWR sky130_fd_sc_hd__decap_12
X_5940_ _5929_/X _5940_/B _5940_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_111_1261 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_890 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1166 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_373 VGND VPWR sky130_fd_sc_hd__decap_12
X_5871_ _5863_/X _5864_/X _5863_/X _5864_/X _5871_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_209_1034 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_905 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_562 VGND VPWR sky130_fd_sc_hd__decap_12
X_7610_ _7227_/X _7160_/A _7729_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4822_ _4822_/A _4821_/X _4887_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_7541_ _7541_/HI la_data_out[68] VGND VPWR sky130_fd_sc_hd__conb_1
X_4753_ _4740_/X _4746_/X _4740_/X _4746_/X _4753_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_187_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_314 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_971 VGND VPWR sky130_fd_sc_hd__decap_12
X_3704_ wbs_adr_i[24] wbs_adr_i[27] wbs_adr_i[26] wbs_adr_i[29] _3704_/X VGND VPWR
+ sky130_fd_sc_hd__or4_4
X_7472_ _7472_/HI io_out[37] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_179_1111 VGND VPWR sky130_fd_sc_hd__decap_6
X_4684_ _4589_/X _4593_/X _4589_/X _4593_/X _4684_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_190_902 VGND VPWR sky130_fd_sc_hd__decap_12
X_6423_ _7714_/Q la_data_in[112] _6487_/A VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_146_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_6354_ _6354_/A _6352_/X _6353_/Y _6354_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_161_147 VGND VPWR sky130_fd_sc_hd__decap_12
X_5305_ _5303_/X _5304_/X _5532_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_142_361 VGND VPWR sky130_fd_sc_hd__decap_12
X_6285_ _5909_/X _5986_/X _5909_/X _5986_/X _6285_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_143_895 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_115_586 VGND VPWR sky130_fd_sc_hd__decap_12
X_5236_ _5233_/X _5234_/X _5235_/X _5236_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_88_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1060 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_1180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_971 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1274 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_1093 VGND VPWR sky130_fd_sc_hd__decap_4
X_5167_ _5160_/X _5166_/X _5160_/X _5166_/X _5167_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_1112 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1127 VGND VPWR sky130_fd_sc_hd__decap_12
X_4118_ _4114_/X _4116_/X _4117_/X _4118_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_5098_ _5093_/X _5097_/X _5093_/X _5097_/X _5098_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_84_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_356 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_507 VGND VPWR sky130_fd_sc_hd__decap_12
X_4049_ _4609_/A _4122_/B _4049_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_72_849 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_501 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_204 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_916 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_215 VGND VPWR sky130_fd_sc_hd__decap_3
X_7808_ _3791_/Y _7808_/Q _7806_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_226 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_409 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_269 VGND VPWR sky130_fd_sc_hd__decap_12
X_7739_ _6350_/Y _4143_/A _7806_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_12_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_612 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_1064 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_166_943 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_870 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_603 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_486 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1217 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_648 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_135 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_564 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_501 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1250 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_971 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_875 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1144 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1166 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_857 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_323 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_627 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_1136 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_367 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_518 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_702 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_556 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_877 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_80 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1202 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_960 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_1008 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_818 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1150 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_1041 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_990 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_681 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1036 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_6070_ _6070_/A _6317_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_190 VGND VPWR sky130_fd_sc_hd__decap_8
X_5021_ _4955_/X _4960_/X _4954_/X _4961_/X _5021_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_100_729 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_418 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_621 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_1217 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_805 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_315 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_529 VGND VPWR sky130_fd_sc_hd__decap_12
X_6972_ _6959_/Y _6960_/Y _6961_/X _6971_/X _7021_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_54_849 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1020 VGND VPWR sky130_fd_sc_hd__decap_6
X_5923_ _5897_/X _5900_/X _5901_/X _5923_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_181_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1121 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_1064 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1079 VGND VPWR sky130_fd_sc_hd__decap_6
X_5854_ _5823_/X _5852_/X _5823_/X _5852_/X _5854_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_146_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_814 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_825 VGND VPWR sky130_fd_sc_hd__decap_3
X_4805_ _4736_/X _4802_/X _4803_/X _4804_/X _4806_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_21_245 VGND VPWR sky130_fd_sc_hd__decap_12
X_5785_ _5730_/X _5734_/X _5730_/X _5734_/X _5785_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_181_1089 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_943 VGND VPWR sky130_fd_sc_hd__decap_3
X_7524_ _7524_/HI la_data_out[51] VGND VPWR sky130_fd_sc_hd__conb_1
X_4736_ _4731_/X _4732_/X _4731_/X _4732_/X _4736_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_175_740 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_289 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_464 VGND VPWR sky130_fd_sc_hd__decap_12
X_7455_ _7455_/HI io_out[20] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_107_306 VGND VPWR sky130_fd_sc_hd__decap_12
X_4667_ _4667_/A _4657_/B _4667_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_119_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_163_946 VGND VPWR sky130_fd_sc_hd__decap_12
X_6406_ _7720_/Q _6408_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_162_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_743 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_659 VGND VPWR sky130_fd_sc_hd__decap_12
X_7386_ io_in[31] _7386_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4598_ _4596_/X _4597_/X _4598_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_150_618 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1122 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_192_1130 VGND VPWR sky130_fd_sc_hd__decap_8
X_6337_ _4123_/B _6334_/B _6337_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_66_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1245 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_89_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_1128 VGND VPWR sky130_fd_sc_hd__decap_8
X_6268_ _6219_/X _6266_/X _6267_/X _7758_/D VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_153_1147 VGND VPWR sky130_fd_sc_hd__decap_12
X_5219_ _5214_/X _5217_/X _5214_/X _5217_/X _5219_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6199_ _6010_/B _6198_/X _6199_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_28_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_996 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_337 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1246 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_724 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_1216 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_554 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_869 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_902 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_784 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_934 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_197_1074 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1121 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1069 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_670 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_488 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_865 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_342 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_171_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_683 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_790 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_900 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_974 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_101 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_1048 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_432 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_668 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_882 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_90_498 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_239 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_598 VGND VPWR sky130_fd_sc_hd__decap_12
X_5570_ _5567_/X _5568_/X _5567_/X _5568_/X _5570_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_79_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_141_1062 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_464 VGND VPWR sky130_fd_sc_hd__decap_12
X_4521_ _4518_/X _4519_/X _4538_/A _4521_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_145_924 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_626 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_783 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_434 VGND VPWR sky130_fd_sc_hd__decap_12
X_7240_ _7187_/X _7239_/X _6085_/X _7240_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_171_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_968 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_1008 VGND VPWR sky130_fd_sc_hd__fill_1
X_4452_ _4653_/A _4546_/B _4452_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_7_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_629 VGND VPWR sky130_fd_sc_hd__decap_12
X_7171_ _7169_/Y _7170_/Y _7169_/Y _7170_/Y _7235_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_4383_ _4323_/X _4381_/X _4378_/X _4382_/X _4383_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_113_843 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_532 VGND VPWR sky130_fd_sc_hd__decap_4
X_6122_ _6089_/X _6120_/X _6121_/X _7782_/D VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_140_662 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_876 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_887 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_576 VGND VPWR sky130_fd_sc_hd__decap_4
X_6053_ _3909_/Y _6058_/B _6053_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_105_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1150 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1233 VGND VPWR sky130_fd_sc_hd__decap_12
X_5004_ _4997_/X _4998_/X _4996_/X _4999_/X _5005_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_152_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_142 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_996 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1186 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_484 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_944 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_148_1216 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_980 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_27 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6955_ _6953_/Y _6954_/Y _6953_/Y _6954_/Y _6955_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_3519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_1129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_476 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_318 VGND VPWR sky130_fd_sc_hd__decap_3
X_5906_ _5885_/X _5905_/X _5885_/X _5905_/X _5906_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_2818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6886_ _6821_/X _6880_/B _6886_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XPHY_2829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_532 VGND VPWR sky130_fd_sc_hd__decap_8
X_5837_ _5834_/X _5835_/X _5836_/X _5837_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_194_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_727 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_666 VGND VPWR sky130_fd_sc_hd__decap_12
X_5768_ _5510_/X _5511_/X _5510_/X _5511_/X _5768_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_136_902 VGND VPWR sky130_fd_sc_hd__fill_1
X_7507_ _7507_/HI la_data_out[34] VGND VPWR sky130_fd_sc_hd__conb_1
X_4719_ _4717_/X _4718_/X _4719_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_5_208 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_795 VGND VPWR sky130_fd_sc_hd__decap_8
X_5699_ _5697_/X _5699_/B _5699_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_108_637 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_1203 VGND VPWR sky130_fd_sc_hd__decap_12
X_7438_ io_oeb[33] _7438_/LO VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_107_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_810 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_403 VGND VPWR sky130_fd_sc_hd__decap_8
X_7369_ _5292_/Y _7355_/X _7368_/X wbs_dat_o[19] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_146_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_990 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_414 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_876 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_342 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_407 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1075 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1086 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1250 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_440 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_760 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_473 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_101 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_175 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_43 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_635 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_977 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_4743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_605 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_487 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_329 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_510 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_4787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_830 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_543 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_201_644 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_200_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_507 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_367 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_199_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_762 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1265 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_570 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_798 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1025 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_802 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_727 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_513 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_1028 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_846 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_922 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_777 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_243 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_741 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_443 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1091 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_178 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_318 VGND VPWR sky130_fd_sc_hd__decap_4
X_6740_ la_data_in[36] _6740_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_3952_ _3951_/A _3951_/B _3951_/X _3952_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_182_1151 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_204_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_684 VGND VPWR sky130_fd_sc_hd__decap_8
X_6671_ _6659_/X _6669_/X _6670_/X _6671_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_3883_ wbs_dat_i[3] _3882_/X _3884_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_176_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1187 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_351 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_1198 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1089 VGND VPWR sky130_fd_sc_hd__decap_8
X_5622_ _4666_/A _5300_/B _5622_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_143_1179 VGND VPWR sky130_fd_sc_hd__decap_12
X_5553_ _5322_/X _5323_/X _5313_/X _5324_/X _5553_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_145_710 VGND VPWR sky130_fd_sc_hd__decap_12
X_4504_ _4499_/A _4498_/B _4506_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_145_754 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_979 VGND VPWR sky130_fd_sc_hd__fill_2
X_5484_ _5483_/A _5482_/X _5483_/X _5484_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_133_916 VGND VPWR sky130_fd_sc_hd__decap_12
X_7223_ _7198_/X _7221_/X _7222_/Y _7612_/D VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_117_489 VGND VPWR sky130_fd_sc_hd__decap_12
X_4435_ _4418_/X _4419_/X _4420_/X _4430_/X _4436_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_104_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_7154_ _7154_/A _7154_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_154_1231 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1234 VGND VPWR sky130_fd_sc_hd__decap_12
X_4366_ _4959_/A _4366_/B _4366_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_6105_ _6100_/X _6102_/Y _6104_/X _7785_/D VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_154_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_215 VGND VPWR sky130_fd_sc_hd__decap_8
X_7085_ _7058_/Y _7060_/B _7060_/X _7084_/X _7085_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_4297_ _4901_/A _4613_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_6036_ _6036_/A _3700_/X _3707_/X _7264_/A VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_86_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1051 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_977 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_13 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_35 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_178 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_46 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_947 VGND VPWR sky130_fd_sc_hd__decap_12
X_6938_ _7644_/Q _6940_/A VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_57 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_68 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_79 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_852 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_931 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_159 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6869_ _6846_/Y _6847_/Y _6868_/X _6869_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XPHY_1914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_323 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_210_430 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1257 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_986 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_1219 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_395 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_474 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_195_698 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_890 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1025 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_746 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_104_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_767 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_778 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_395 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_922 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_703 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_635 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_741 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_251 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_487 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_960 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_446 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_993 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_621 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_492 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_975 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1029 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1062 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1182 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_1242 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_787 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_177_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1158 VGND VPWR sky130_fd_sc_hd__decap_12
X_4220_ _4219_/A _4219_/B _4219_/X _4220_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_141_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_159 VGND VPWR sky130_fd_sc_hd__decap_12
X_4151_ _4110_/X _4149_/X _4110_/X _4149_/X _4151_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_96_833 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_877 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_568 VGND VPWR sky130_fd_sc_hd__decap_12
X_4082_ _4793_/A _4123_/B _4082_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_62_1180 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_1153 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_110_1123 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_955 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1247 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_1227 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_184_1235 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_947 VGND VPWR sky130_fd_sc_hd__decap_12
X_7772_ _7772_/D _4886_/A _7774_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_145_1219 VGND VPWR sky130_fd_sc_hd__fill_1
X_4984_ _4943_/X _4944_/X _4943_/X _4944_/X _4986_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6723_ _6723_/A _6723_/B _6723_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_3935_ _3927_/X _3926_/X _3934_/X _3935_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_211_249 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_345 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1063 VGND VPWR sky130_fd_sc_hd__decap_4
X_6654_ _6618_/Y _6619_/Y _6685_/B _6654_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_3866_ _6333_/A _3866_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_5605_ _5480_/X _5484_/X _5480_/X _5484_/X _5605_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6585_ _6521_/X _6541_/B _6585_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
X_3797_ _3757_/A _3798_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_164_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_220 VGND VPWR sky130_fd_sc_hd__decap_12
X_5536_ _5532_/X _5533_/X _5534_/Y _5535_/X _5536_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_133_702 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_724 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_938 VGND VPWR sky130_fd_sc_hd__decap_8
X_5467_ _5233_/A _4844_/B _5467_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_105_426 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_160_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_757 VGND VPWR sky130_fd_sc_hd__decap_12
X_7206_ la_data_in[111] _7207_/B _7206_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_4418_ _4412_/X _4413_/X _4411_/X _4414_/X _4418_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_5398_ _6228_/A _6223_/A _6008_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_114_971 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_513 VGND VPWR sky130_fd_sc_hd__decap_3
X_7137_ _6052_/A _7210_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_113_470 VGND VPWR sky130_fd_sc_hd__decap_12
X_4349_ _4280_/X _4281_/X _4280_/X _4281_/X _4349_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_87_855 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_643 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_708 VGND VPWR sky130_fd_sc_hd__decap_12
X_7068_ la_data_in[83] _7068_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_6019_ _6019_/A _6019_/B _6019_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_86_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_56 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_605 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_3102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_28_999 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_722 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_245 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_593 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_788 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_146_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1024 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_991 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_440 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_44 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_507 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_304 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_315 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1040 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_837 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_398 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_182_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_690 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_757 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1022 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_597 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_9 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_1028 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_538 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_571 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_733 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_276 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_643 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1252 VGND VPWR sky130_fd_sc_hd__decap_12
X_3720_ _3720_/A _4565_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_187_963 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_163 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_123 VGND VPWR sky130_fd_sc_hd__decap_12
X_6370_ _4959_/B _6373_/B _6372_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_61_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_871 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_562 VGND VPWR sky130_fd_sc_hd__decap_12
X_5321_ _5319_/X _5320_/X _5319_/X _5320_/X _5321_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_177_1050 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_852 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_391 VGND VPWR sky130_fd_sc_hd__decap_12
X_5252_ _5108_/X _5112_/X _5108_/X _5112_/X _5252_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_170_896 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_727 VGND VPWR sky130_fd_sc_hd__decap_12
X_4203_ _4069_/X _4096_/X _4104_/A _4203_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_190_1250 VGND VPWR sky130_fd_sc_hd__fill_1
X_5183_ _5174_/X _5182_/X _5174_/X _5182_/X _5183_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_151_1212 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_630 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_855 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_708 VGND VPWR sky130_fd_sc_hd__decap_12
X_4134_ _4841_/A _4277_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_888 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_825 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_313 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_847 VGND VPWR sky130_fd_sc_hd__decap_12
X_4065_ _4039_/X _4064_/X _4065_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_113_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1130 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_251 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_593 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_284 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_1095 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_408 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_969 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_51_232 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_419 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_149_1196 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_608 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_788 VGND VPWR sky130_fd_sc_hd__decap_12
X_4967_ _4963_/X _4966_/X _4963_/X _4966_/X _4967_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7755_ _7755_/D _5751_/A _7754_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_1213 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3918_ _4189_/A _3918_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_6706_ _6694_/X _6643_/X _6705_/Y _6706_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_7686_ _7686_/D _6630_/A _7658_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4898_ _4898_/A _4959_/B _4824_/A _4898_/D _4949_/B VGND VPWR sky130_fd_sc_hd__or4_4
X_6637_ la_data_in[18] _6638_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_165_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_410 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_849 VGND VPWR sky130_fd_sc_hd__decap_12
X_3849_ _3832_/A _3847_/X _3849_/C _3849_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_193_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_819 VGND VPWR sky130_fd_sc_hd__decap_12
X_6568_ _6501_/A la_data_in[11] _6503_/X _6568_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_146_860 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1131 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_306 VGND VPWR sky130_fd_sc_hd__decap_12
X_5519_ _5516_/A _5516_/B _5518_/Y _6198_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_161_830 VGND VPWR sky130_fd_sc_hd__decap_12
X_6499_ la_data_in[12] _6500_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_195_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_373 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_730 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_880 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_571 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_716 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_525 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_87 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_569 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_939 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_449 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_27 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_922 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_601 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_623 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_337 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_627 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_1128 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1248 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_727 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_873 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_803 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_611 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_516 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1101 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_730 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_508 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_251 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_1273 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_1224 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1178 VGND VPWR sky130_fd_sc_hd__decap_12
X_5870_ _5827_/X _5828_/X _5829_/X _5870_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_80_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_917 VGND VPWR sky130_fd_sc_hd__decap_4
X_4821_ _4821_/A _5301_/B _4821_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_178_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_574 VGND VPWR sky130_fd_sc_hd__decap_12
X_7540_ _7540_/HI la_data_out[67] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_159_440 VGND VPWR sky130_fd_sc_hd__decap_8
X_4752_ _4747_/X _4751_/X _4747_/X _4751_/X _4752_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_119_304 VGND VPWR sky130_fd_sc_hd__fill_1
X_3703_ wbs_adr_i[28] wbs_adr_i[31] _3706_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_174_410 VGND VPWR sky130_fd_sc_hd__decap_12
X_7471_ _7471_/HI io_out[36] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_105_1044 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_983 VGND VPWR sky130_fd_sc_hd__decap_12
X_4683_ _4678_/X _4682_/X _4681_/X _4683_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_6422_ la_data_in[113] _6422_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_175_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_914 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1099 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_638 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_190_947 VGND VPWR sky130_fd_sc_hd__decap_12
X_6353_ wbs_dat_i[8] _6349_/B _6353_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_162_649 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_830 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_841 VGND VPWR sky130_fd_sc_hd__decap_12
X_5304_ _5304_/A _4492_/A _5304_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_161_159 VGND VPWR sky130_fd_sc_hd__decap_12
X_6284_ _6282_/Y _6283_/X _7755_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_130_502 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_5235_ _5233_/X _5234_/X _5235_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_9_1253 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_579 VGND VPWR sky130_fd_sc_hd__fill_1
X_5166_ _5161_/X _5165_/X _5161_/X _5165_/X _5166_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_5_1117 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_1124 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_1139 VGND VPWR sky130_fd_sc_hd__decap_12
X_4117_ _4114_/X _4116_/X _4117_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_83_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1037 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_335 VGND VPWR sky130_fd_sc_hd__fill_1
X_5097_ _5096_/A _5096_/B _5096_/X _5097_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_186_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_666 VGND VPWR sky130_fd_sc_hd__decap_12
X_4048_ _4041_/X _4047_/X _4041_/X _4047_/X _4048_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_204_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_58 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_861 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_216 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_703 VGND VPWR sky130_fd_sc_hd__decap_12
X_7807_ _3801_/Y _7807_/Q _7806_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_227 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_928 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_546 VGND VPWR sky130_fd_sc_hd__decap_3
X_5999_ _5993_/X _5998_/Y _6000_/D VGND VPWR sky130_fd_sc_hd__and2_4
XPHY_238 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_276 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_249 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_1130 VGND VPWR sky130_fd_sc_hd__decap_12
X_7738_ _6354_/Y _7738_/Q _7806_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_166_911 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_281 VGND VPWR sky130_fd_sc_hd__decap_12
X_7669_ _6808_/X _6742_/A _7707_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_137_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_914 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_679 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_1188 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_999 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_192_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_318 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_615 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1229 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_690 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_109_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_532 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_340 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_405 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_682 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_43 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_803 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1123 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_983 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_887 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1156 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_335 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_869 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_349 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_541 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1044 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_574 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_568 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_771 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_602 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1090 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_1214 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_910 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_972 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_292 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_1138 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_977 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_209_27 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_102_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_785 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1001 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1020 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_143_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_703 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1053 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_693 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_257 VGND VPWR sky130_fd_sc_hd__decap_12
X_5020_ _7774_/Q _5020_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_112_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_817 VGND VPWR sky130_fd_sc_hd__decap_6
X_6971_ _6962_/Y _6963_/Y _6964_/X _6970_/X _6971_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_53_327 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_647 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_891 VGND VPWR sky130_fd_sc_hd__decap_12
X_5922_ _5918_/X _5919_/X _5920_/Y _5921_/X _5922_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_207_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_390 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_185_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1013 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1185 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_703 VGND VPWR sky130_fd_sc_hd__decap_12
X_5853_ _5839_/X _5848_/X _5847_/X _5849_/X _5853_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_107_1106 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_1166 VGND VPWR sky130_fd_sc_hd__fill_1
X_4804_ _4736_/X _4802_/X _4736_/X _4802_/X _4804_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_142_1008 VGND VPWR sky130_fd_sc_hd__decap_12
X_5784_ _5742_/X _5743_/X _5742_/X _5743_/X _5784_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_148_911 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_257 VGND VPWR sky130_fd_sc_hd__fill_1
X_4735_ _4544_/X _4734_/X _4544_/X _4734_/X _4806_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7523_ _7523_/HI la_data_out[50] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_159_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_752 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_808 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_27 VGND VPWR sky130_fd_sc_hd__decap_12
X_7454_ _7454_/HI io_out[19] VGND VPWR sky130_fd_sc_hd__conb_1
X_4666_ _4666_/A _4666_/B _4666_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_174_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_318 VGND VPWR sky130_fd_sc_hd__decap_12
X_6405_ _6403_/Y _6405_/B _6405_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_163_958 VGND VPWR sky130_fd_sc_hd__decap_12
X_7385_ _4580_/Y _7354_/X _7384_/X wbs_dat_o[24] VGND VPWR sky130_fd_sc_hd__o21ai_4
X_4597_ _4514_/A _4597_/B _4597_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_162_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_755 VGND VPWR sky130_fd_sc_hd__decap_8
X_6336_ _6350_/A _6336_/B _6335_/Y _6336_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_143_660 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_202 VGND VPWR sky130_fd_sc_hd__decap_12
X_6267_ _5632_/Y _6216_/X _6194_/X _6267_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_115_395 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_855 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_557 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_877 VGND VPWR sky130_fd_sc_hd__decap_12
X_5218_ _5072_/X _5076_/X _5072_/X _5076_/X _5218_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6198_ _6198_/A _6198_/B _6008_/A _6197_/X _6198_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_57_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_398 VGND VPWR sky130_fd_sc_hd__decap_12
X_5149_ _5078_/X _5082_/X _5081_/X _5149_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_84_430 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_666 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_880 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_1230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_530 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1116 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_56 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_680 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_78 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_566 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_538 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_944 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_914 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_711 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_627 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_682 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_833 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_912 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_986 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_989 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_833 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_574 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1249 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_188_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_196 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_870 VGND VPWR sky130_fd_sc_hd__decap_12
X_4520_ _4518_/X _4519_/X _4538_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_8_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_156_251 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1074 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_638 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1099 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_593 VGND VPWR sky130_fd_sc_hd__decap_12
X_4451_ _4386_/X _4441_/X _4444_/Y _4451_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_102_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_232 VGND VPWR sky130_fd_sc_hd__decap_12
X_7170_ la_data_in[101] _7170_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_113_800 VGND VPWR sky130_fd_sc_hd__fill_1
X_4382_ _4323_/X _4381_/X _4323_/X _4381_/X _4382_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_98_500 VGND VPWR sky130_fd_sc_hd__fill_1
X_6121_ _4070_/Y _6103_/X _6092_/X _6121_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_113_855 VGND VPWR sky130_fd_sc_hd__decap_12
X_6052_ _6052_/A _6057_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_100_505 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_588 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_899 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_739 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_611 VGND VPWR sky130_fd_sc_hd__decap_12
X_5003_ _7775_/Q _5003_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_112_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1162 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1245 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_1109 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_305 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1198 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_496 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_293 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1228 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_658 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_349 VGND VPWR sky130_fd_sc_hd__decap_12
X_6954_ la_data_in[69] _6954_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_208_992 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_5905_ _5886_/X _5904_/X _5905_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_2808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6885_ _6885_/A _6883_/Y _6885_/C _7665_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_179_354 VGND VPWR sky130_fd_sc_hd__decap_12
X_5836_ _5834_/X _5835_/X _5836_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_61_190 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_324 VGND VPWR sky130_fd_sc_hd__decap_12
X_5767_ _5513_/X _5514_/X _5513_/X _5514_/X _5767_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_10_739 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_678 VGND VPWR sky130_fd_sc_hd__decap_12
X_7506_ _7506_/HI la_data_out[33] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_108_605 VGND VPWR sky130_fd_sc_hd__decap_12
X_4718_ _4718_/A _4743_/B _4718_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_5698_ _5216_/A _4595_/B _5699_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_163_733 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_194_1215 VGND VPWR sky130_fd_sc_hd__decap_12
X_4649_ _4655_/A _4657_/B _4649_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7437_ io_oeb[32] _7437_/LO VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_107_159 VGND VPWR sky130_fd_sc_hd__decap_12
X_7368_ _5294_/A _7349_/X _7367_/Y _7364_/X _7368_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_162_276 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_426 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1070 VGND VPWR sky130_fd_sc_hd__fill_1
X_6319_ _6319_/A _7730_/Q _6319_/C _7746_/Q _6319_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_7299_ io_in[12] _7299_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_131_641 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_685 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_1115 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_975 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1137 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_772 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_154 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_176_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_485 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_33 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_422 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_55 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_45_647 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_444 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_428 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_617 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1071 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1044 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_1172 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_623 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_190 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_515 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_656 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1260 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1233 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_774 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_936 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_593 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1012 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_972 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_814 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_971 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_1059 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_858 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_750 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_233 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_255 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_934 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_789 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_455 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_1160 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_263 VGND VPWR sky130_fd_sc_hd__decap_12
X_3951_ _3951_/A _3951_/B _3951_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_189_663 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_138 VGND VPWR sky130_fd_sc_hd__decap_12
X_6670_ _6670_/A _6670_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_91_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_3882_ _3759_/A _3882_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_204_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_886 VGND VPWR sky130_fd_sc_hd__decap_12
X_5621_ _4667_/A _5301_/B _5623_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_176_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_363 VGND VPWR sky130_fd_sc_hd__decap_3
X_5552_ _5529_/X _5530_/X _5529_/X _5530_/X _5552_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_145_722 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_582 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_947 VGND VPWR sky130_fd_sc_hd__decap_12
X_4503_ _4503_/A _4497_/B _4503_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_145_733 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_581 VGND VPWR sky130_fd_sc_hd__decap_12
X_5483_ _5483_/A _5482_/X _5483_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_145_766 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_457 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_703 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_928 VGND VPWR sky130_fd_sc_hd__decap_8
X_4434_ _4434_/A _4434_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_7222_ _7198_/X _7221_/X _7212_/X _7222_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_144_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_7153_ _7151_/Y _7152_/Y _7153_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_4365_ _4497_/B _4366_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_154_1243 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_1246 VGND VPWR sky130_fd_sc_hd__decap_4
X_6104_ _3988_/Y _6103_/X _6092_/X _6104_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_7084_ _7061_/Y _7062_/Y _7083_/X _7084_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_4296_ _4295_/Y _4901_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_154_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_836 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1020 VGND VPWR sky130_fd_sc_hd__decap_12
X_6035_ wbs_adr_i[4] _6036_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_55_901 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_794 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_731 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_1063 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_26_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_764 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_14 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_989 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_25 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_36 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6937_ _6935_/Y _6937_/B _6937_/X VGND VPWR sky130_fd_sc_hd__and2_4
XPHY_2605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_148_1069 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_820 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_959 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_69 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_611 VGND VPWR sky130_fd_sc_hd__decap_8
X_6868_ _6911_/A _6867_/X _6868_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_1915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_943 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_184 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_442 VGND VPWR sky130_fd_sc_hd__decap_12
X_5819_ _5781_/X _5817_/X _5819_/X VGND VPWR sky130_fd_sc_hd__and2_4
XPHY_1948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_806 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_694 VGND VPWR sky130_fd_sc_hd__decap_8
X_6799_ _7672_/Q la_data_in[38] _6735_/X _6799_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_194_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_379 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_183_828 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_486 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_148_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_958 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1034 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1037 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1089 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_758 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_245 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_983 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_674 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_696 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1062 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_934 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_591 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_444 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_263 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_105 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_948 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_269 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_972 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_4596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_330 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_471 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_633 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_987 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_891 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_139_582 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1191 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1074 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_142_703 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1254 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_265 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_276 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_747 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_257 VGND VPWR sky130_fd_sc_hd__decap_12
X_4150_ _7781_/Q _4150_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_122_471 VGND VPWR sky130_fd_sc_hd__decap_12
X_4081_ _4539_/A _4122_/B _4081_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_55_208 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_271 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_586 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_967 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1259 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_184_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_753 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_403 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_617 VGND VPWR sky130_fd_sc_hd__decap_12
X_7771_ _7771_/D _4812_/A _7774_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_36_499 VGND VPWR sky130_fd_sc_hd__fill_1
X_4983_ _6015_/A _4982_/X _4983_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_52_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_138 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_781 VGND VPWR sky130_fd_sc_hd__decap_12
X_6722_ la_data_in[42] _6723_/B VGND VPWR sky130_fd_sc_hd__inv_8
X_3934_ _3722_/A _3949_/B _4609_/A _3933_/X _3934_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_32_650 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_823 VGND VPWR sky130_fd_sc_hd__fill_1
X_3865_ _3832_/A _3865_/B _3865_/C _7799_/D VGND VPWR sky130_fd_sc_hd__nor3_4
X_6653_ _6620_/X _6684_/B _6685_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_32_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_149_357 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_176_154 VGND VPWR sky130_fd_sc_hd__decap_12
X_5604_ _5601_/X _5602_/X _5603_/X _5604_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_20_867 VGND VPWR sky130_fd_sc_hd__decap_12
X_3796_ _5052_/A _4467_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_6584_ _6542_/X _6582_/X _6583_/Y _6584_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_164_349 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_191_135 VGND VPWR sky130_fd_sc_hd__decap_12
X_5535_ _5532_/X _5533_/X _5532_/X _5533_/X _5535_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_145_541 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_788 VGND VPWR sky130_fd_sc_hd__decap_8
X_5466_ _5176_/A _4847_/B _5466_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_132_202 VGND VPWR sky130_fd_sc_hd__decap_12
X_4417_ _4390_/X _4405_/X _4415_/X _4416_/X _4417_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_7205_ io_out[6] _7204_/X _7207_/B VGND VPWR sky130_fd_sc_hd__xnor2_4
XFILLER_160_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_769 VGND VPWR sky130_fd_sc_hd__decap_12
X_5397_ _6005_/A _6005_/B _5396_/Y _6223_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_120_419 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1160 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_672 VGND VPWR sky130_fd_sc_hd__decap_12
X_4348_ _4337_/X _4338_/X _4336_/X _4348_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_7136_ _7078_/X _7134_/X _7135_/Y _7620_/D VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_143_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_611 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_8_1137 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_482 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_867 VGND VPWR sky130_fd_sc_hd__decap_12
X_7067_ _7621_/Q _7067_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4279_ _4276_/X _4279_/B _4279_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_143_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_1008 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1019 VGND VPWR sky130_fd_sc_hd__decap_12
X_6018_ _6018_/A _6018_/B _6018_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_55_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_414 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_105 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_734 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_3136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_257 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_408 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1172 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1183 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_661 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_672 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1036 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_193 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_733 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_849 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_755 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_308 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_703 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_170_319 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_510 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_566 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1034 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_780 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_753 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_550 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_556 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_583 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_274 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_745 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_611 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_3670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_655 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_187_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_182 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_828 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_175 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_174_658 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_530 VGND VPWR sky130_fd_sc_hd__decap_12
X_5320_ _5175_/X _5181_/X _5174_/X _5182_/X _5320_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_6_860 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3 VGND VPWR sky130_fd_sc_hd__decap_4
X_5251_ _5231_/X _5239_/X _5249_/X _5250_/X _5251_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_142_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_886 VGND VPWR sky130_fd_sc_hd__decap_3
X_4202_ _4200_/X _4201_/X _4202_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_64_1243 VGND VPWR sky130_fd_sc_hd__decap_8
X_5182_ _5175_/X _5181_/X _5175_/X _5181_/X _5182_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_130_739 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_642 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_1276 VGND VPWR sky130_fd_sc_hd__fill_1
X_4133_ _7738_/Q _4841_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_111_975 VGND VPWR sky130_fd_sc_hd__fill_1
X_4064_ _4040_/X _4061_/X _4062_/X _4063_/X _4064_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_110_485 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_859 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_325 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_1191 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1044 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_409 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_91_391 VGND VPWR sky130_fd_sc_hd__fill_1
X_7754_ _6287_/Y _5807_/A _7754_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4966_ _4964_/X _4965_/X _4964_/X _4965_/X _4966_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_196_227 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1225 VGND VPWR sky130_fd_sc_hd__fill_1
X_6705_ _6705_/A _6642_/X _6705_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_51_288 VGND VPWR sky130_fd_sc_hd__decap_12
X_3917_ _4583_/A _4189_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_7685_ _7685_/D _6633_/A _7658_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4897_ _4609_/A _4959_/B _4959_/A _4898_/D _4897_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_32_491 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_642 VGND VPWR sky130_fd_sc_hd__decap_12
X_6636_ _7684_/Q _6636_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_177_485 VGND VPWR sky130_fd_sc_hd__decap_3
X_3848_ wbs_dat_i[7] _3848_/B _3849_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_138_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1050 VGND VPWR sky130_fd_sc_hd__decap_12
X_3779_ _4513_/A _4769_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_6567_ _6550_/X _6565_/X _6566_/Y _6567_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_193_989 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_4_808 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_552 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_146_872 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_703 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_1_0_wb_clk_i clkbuf_3_0_0_wb_clk_i/X _7707_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_5518_ _5518_/A _5518_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_180_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_318 VGND VPWR sky130_fd_sc_hd__decap_12
X_6498_ _6498_/A _6500_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_173_691 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_190 VGND VPWR sky130_fd_sc_hd__decap_12
X_5449_ _5447_/X _5448_/X _5447_/X _5448_/X _5449_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_105_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_227 VGND VPWR sky130_fd_sc_hd__decap_12
X_7119_ _7119_/A _7119_/B _7120_/C VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_86_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_56 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_1062 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_807 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_742 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_764 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_904 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1242 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_892 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_583 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_723 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_959 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_728 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_537 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_99 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_288 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_761 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_635 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_155_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_349 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_174 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_184_978 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1112 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_196 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1156 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1224 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_907 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_330 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_340 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_1219 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_588 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_351 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_739 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_896 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_815 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_1129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_686 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1113 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_818 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_689 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_1203 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1003 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_1236 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_391 VGND VPWR sky130_fd_sc_hd__decap_3
X_4820_ _4820_/A _4820_/B _4822_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_22_929 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1069 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_586 VGND VPWR sky130_fd_sc_hd__decap_3
X_4751_ _4748_/X _4749_/X _4750_/X _4751_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_105_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_951 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_202_581 VGND VPWR sky130_fd_sc_hd__decap_8
X_3702_ wbs_adr_i[5] wbs_adr_i[7] wbs_adr_i[6] wbs_adr_i[17] _3702_/X VGND VPWR sky130_fd_sc_hd__or4_4
X_4682_ _4679_/X _4680_/X _4681_/X _4682_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_7470_ _7470_/HI io_out[35] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_187_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1094 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_995 VGND VPWR sky130_fd_sc_hd__decap_12
X_6421_ _6421_/A _6421_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_135_809 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_606 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_926 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_488 VGND VPWR sky130_fd_sc_hd__decap_12
X_6352_ _4137_/X _6348_/B _6352_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_190_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_522 VGND VPWR sky130_fd_sc_hd__decap_12
X_5303_ _5300_/X _5301_/X _5532_/A _5303_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_154_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_853 VGND VPWR sky130_fd_sc_hd__fill_1
X_6283_ _5751_/Y _6091_/X _6208_/A _6283_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_130_514 VGND VPWR sky130_fd_sc_hd__decap_4
X_5234_ _5234_/A _4748_/B _5234_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_142_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1130 VGND VPWR sky130_fd_sc_hd__decap_12
X_5165_ _5162_/X _5163_/X _5164_/X _5165_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_111_750 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_141 VGND VPWR sky130_fd_sc_hd__decap_12
X_4116_ _4499_/A _4218_/B _4116_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_111_794 VGND VPWR sky130_fd_sc_hd__decap_12
X_5096_ _5096_/A _5096_/B _5096_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_112_1049 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_15 VGND VPWR sky130_fd_sc_hd__decap_4
X_4047_ _4045_/X _4046_/X _4044_/X _4047_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_84_678 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_26 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_550 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_306 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_140_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_745 VGND VPWR sky130_fd_sc_hd__decap_8
X_7806_ _3809_/Y _7806_/Q _7806_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_206 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_873 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_228 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_715 VGND VPWR sky130_fd_sc_hd__decap_4
X_5998_ _5998_/A _5998_/B _5997_/Y _5998_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XPHY_239 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_507 VGND VPWR sky130_fd_sc_hd__decap_12
X_7737_ _6357_/Y _7737_/Q _7806_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_36_1142 VGND VPWR sky130_fd_sc_hd__decap_12
X_4949_ _4949_/A _4949_/B _5023_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_21_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_923 VGND VPWR sky130_fd_sc_hd__decap_12
X_7668_ _6813_/X _6745_/A _7707_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_177_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1099 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_135 VGND VPWR sky130_fd_sc_hd__decap_12
X_6619_ la_data_in[24] _6619_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_7599_ _7599_/HI la_data_out[126] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_192_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_627 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_104 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_352 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_672 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_417 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_161_694 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1162 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_55 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_750 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_815 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_995 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_837 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_623 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_1127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_196 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_347 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_818 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_380 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_167_1050 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_851 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_203 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_288 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_93 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_901 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_759 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_208 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_783 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_794 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_922 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_282 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_984 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_764 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_669 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_989 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_172_937 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_959 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_498 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_447 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1073 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_1065 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1087 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_973 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_464 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_678 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1151 VGND VPWR sky130_fd_sc_hd__decap_4
X_6970_ _6965_/Y _6966_/Y _6969_/X _6970_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_19_550 VGND VPWR sky130_fd_sc_hd__decap_12
X_5921_ _5918_/X _5919_/X _5918_/X _5919_/X _5921_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_53_339 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1172 VGND VPWR sky130_fd_sc_hd__decap_12
X_5852_ _5841_/X _5842_/X _5850_/X _5851_/X _5852_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_181_1025 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_715 VGND VPWR sky130_fd_sc_hd__decap_12
X_4803_ _4797_/X _4798_/X _4796_/X _4799_/X _4803_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_21_225 VGND VPWR sky130_fd_sc_hd__fill_2
X_5783_ _5697_/X _5699_/B _5699_/X _5783_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_194_506 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_1189 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_236 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_923 VGND VPWR sky130_fd_sc_hd__decap_12
X_7522_ _7522_/HI la_data_out[49] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_9_71 VGND VPWR sky130_fd_sc_hd__decap_12
X_4734_ _4711_/X _4733_/X _4711_/X _4733_/X _4734_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_175_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_967 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_119_135 VGND VPWR sky130_fd_sc_hd__decap_12
X_7453_ _7453_/HI io_out[18] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_175_764 VGND VPWR sky130_fd_sc_hd__decap_12
X_4665_ _4665_/A _4665_/B _4665_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_119_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1050 VGND VPWR sky130_fd_sc_hd__decap_8
X_6404_ la_data_in[119] _6405_/B VGND VPWR sky130_fd_sc_hd__inv_8
X_7384_ _3918_/X _7370_/X _7383_/Y _7265_/X _7384_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_4596_ _4513_/A _4596_/B _4596_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_6335_ wbs_dat_i[13] _6338_/B _6335_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_190_778 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_801 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_27 VGND VPWR sky130_fd_sc_hd__decap_12
X_6266_ _5993_/D _5766_/X _5993_/D _5766_/X _6266_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_5217_ _5215_/X _5216_/X _5217_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_103_569 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_889 VGND VPWR sky130_fd_sc_hd__decap_12
X_6197_ _6000_/D _6197_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_57_623 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_1095 VGND VPWR sky130_fd_sc_hd__decap_3
X_5148_ _5143_/X _5147_/X _5143_/X _5147_/X _5148_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_151_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_442 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_678 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_818 VGND VPWR sky130_fd_sc_hd__decap_12
X_5079_ _4667_/A _4844_/B _5079_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_151_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1242 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_840 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_542 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_1275 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_704 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_1128 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_692 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_708 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_578 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_989 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_926 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_617 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_291 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_403 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_723 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_126_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_691 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_812 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_180_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_897 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_652 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_943 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_998 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1241 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1156 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_892 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_648 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1274 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_391 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_204_621 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_147 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_188_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_467 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_862 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_309 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_845 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_654 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_867 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_176_506 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1050 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_411 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1151 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1045 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_882 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_4450_ _4321_/X _4383_/X _4385_/X _4450_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_145_959 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_172_745 VGND VPWR sky130_fd_sc_hd__decap_12
X_4381_ _4324_/X _4375_/X _4379_/X _4380_/X _4381_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_6120_ _4208_/X _6096_/X _4208_/X _6096_/X _6120_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_112_300 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_631 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_322 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_867 VGND VPWR sky130_fd_sc_hd__fill_2
X_6051_ _6044_/A _6052_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_26_1130 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_517 VGND VPWR sky130_fd_sc_hd__fill_2
X_5002_ _4994_/X _4995_/X _5000_/X _5001_/X _5002_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_113_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_943 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_1174 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_317 VGND VPWR sky130_fd_sc_hd__decap_12
X_6953_ _7639_/Q _6953_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_19_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_147 VGND VPWR sky130_fd_sc_hd__fill_2
X_5904_ _5896_/X _5903_/X _5896_/X _5903_/X _5904_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_2809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_489 VGND VPWR sky130_fd_sc_hd__decap_12
X_6884_ la_data_in[63] _6884_/B _6885_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_34_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_62 VGND VPWR sky130_fd_sc_hd__decap_12
X_5835_ _4697_/A _5835_/B _5835_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_139_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_876 VGND VPWR sky130_fd_sc_hd__decap_8
X_5766_ _5725_/X _5762_/X _5765_/Y _5766_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_7505_ _7505_/HI la_data_out[32] VGND VPWR sky130_fd_sc_hd__conb_1
X_4717_ _4697_/A _4666_/B _4717_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_120_1104 VGND VPWR sky130_fd_sc_hd__decap_12
X_5697_ _5215_/A _4137_/X _5697_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_135_403 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_617 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_7436_ io_oeb[31] _7436_/LO VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_190_520 VGND VPWR sky130_fd_sc_hd__decap_12
X_4648_ _4648_/A _4657_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_194_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_929 VGND VPWR sky130_fd_sc_hd__decap_8
X_7367_ io_in[25] _7367_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4579_ _4560_/X _4576_/X _4577_/X _4578_/X _4579_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_89_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_683 VGND VPWR sky130_fd_sc_hd__decap_12
X_6318_ _6316_/Y _6317_/X _6320_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_115_171 VGND VPWR sky130_fd_sc_hd__decap_12
X_7298_ _7784_/Q _7292_/B _7298_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_130_141 VGND VPWR sky130_fd_sc_hd__decap_12
X_6249_ _5779_/X _6248_/X _6249_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_104_889 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_1230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_697 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_987 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_1149 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_784 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_924 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_4701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_946 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_4712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_434 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_659 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_456 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_4745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_1050 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_629 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_1083 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1151 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_331 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_186_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_527 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_668 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_200_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_892 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_414 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_734 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_650 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_298 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1024 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_707 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1098 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_984 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_1008 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_686 VGND VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_14_0_wb_clk_i clkbuf_3_7_0_wb_clk_i/X _7810_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_95_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_757 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_401 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_412 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_114 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_467 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_873 VGND VPWR sky130_fd_sc_hd__decap_12
X_3950_ _4565_/A _3950_/B _3951_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_205_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_361 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1036 VGND VPWR sky130_fd_sc_hd__fill_1
X_3881_ _5185_/A _3897_/B _3884_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_177_826 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1069 VGND VPWR sky130_fd_sc_hd__decap_12
X_5620_ _5615_/X _5619_/X _5618_/X _5620_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_32_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_5551_ _5540_/X _5541_/X _5540_/X _5541_/X _5551_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_157_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_690 VGND VPWR sky130_fd_sc_hd__decap_12
X_4502_ _4497_/X _4501_/X _4497_/X _4501_/X _4502_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_172_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_959 VGND VPWR sky130_fd_sc_hd__decap_12
X_5482_ _4716_/A _4299_/X _5482_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_8_593 VGND VPWR sky130_fd_sc_hd__decap_12
X_7221_ _7154_/A la_data_in[106] _7156_/X _7221_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_117_469 VGND VPWR sky130_fd_sc_hd__decap_12
X_4433_ _4389_/X _4417_/X _4431_/X _4432_/X _4433_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_99_810 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_288 VGND VPWR sky130_fd_sc_hd__fill_2
X_7152_ la_data_in[107] _7152_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4364_ _4612_/B _4497_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_141_940 VGND VPWR sky130_fd_sc_hd__decap_12
X_6103_ _6158_/A _6103_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_140_450 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1258 VGND VPWR sky130_fd_sc_hd__fill_1
X_4295_ _4295_/A _4295_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_7083_ _7083_/A _7083_/B _7083_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_141_984 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_848 VGND VPWR sky130_fd_sc_hd__decap_6
X_6034_ _7327_/A _6034_/B _6034_/C _6034_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_6_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_581 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_743 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_125 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_220 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_15 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_147 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_26 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_199_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_776 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6936_ la_data_in[75] _6937_/B VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_37 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_48 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_681 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_900 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_832 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6867_ _6849_/Y _6850_/Y _6866_/X _6867_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XPHY_2639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_210_410 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1237 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_955 VGND VPWR sky130_fd_sc_hd__decap_6
X_5818_ _5781_/X _5817_/X _5820_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XPHY_1938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_196 VGND VPWR sky130_fd_sc_hd__decap_12
X_6798_ _6760_/X _6796_/X _6797_/Y _6798_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XPHY_1949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_454 VGND VPWR sky130_fd_sc_hd__decap_4
X_5749_ _5749_/A _5749_/B _5749_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_194_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_498 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_414 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_948 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_159_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1240 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_918 VGND VPWR sky130_fd_sc_hd__decap_8
X_7419_ io_oeb[14] _7419_/LO VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_124_929 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1049 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_586 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_1199 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_450 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_995 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_483 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_537 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_434 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_1104 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_456 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_916 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_32 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_489 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_117 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_990 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_459 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_342 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_999 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_201_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_509 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_186_678 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_306 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_701 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_594 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_745 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_759 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_123_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_984 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_483 VGND VPWR sky130_fd_sc_hd__decap_12
X_4080_ _4073_/X _4079_/X _4073_/X _4079_/X _4080_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_1_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_1111 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_510 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_710 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1227 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_581 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_1245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_231 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_776 VGND VPWR sky130_fd_sc_hd__decap_8
X_7770_ _7770_/D _4580_/A _7774_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_24_629 VGND VPWR sky130_fd_sc_hd__decap_12
X_4982_ _4982_/A _4982_/B _4982_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_184_1259 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_670 VGND VPWR sky130_fd_sc_hd__fill_1
X_6721_ _7676_/Q _6723_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_211_218 VGND VPWR sky130_fd_sc_hd__decap_12
X_3933_ _3950_/B _3933_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_6652_ _6621_/Y _6623_/B _6623_/X _6651_/X _6684_/B VGND VPWR sky130_fd_sc_hd__o22a_4
X_3864_ wbs_dat_i[5] _3848_/B _3865_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_60_993 VGND VPWR sky130_fd_sc_hd__decap_12
X_5603_ _5601_/X _5602_/X _5603_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_6583_ _6542_/X _6582_/X _6572_/X _6583_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_176_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_879 VGND VPWR sky130_fd_sc_hd__decap_6
X_3795_ _4554_/A _5052_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_178_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1221 VGND VPWR sky130_fd_sc_hd__decap_12
X_5534_ _5534_/A _5534_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_191_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_406 VGND VPWR sky130_fd_sc_hd__decap_12
X_5465_ _5408_/X _5412_/X _5408_/X _5412_/X _5465_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_172_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_428 VGND VPWR sky130_fd_sc_hd__decap_12
X_7204_ _7142_/Y _7143_/Y _7203_/X _7204_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_4416_ _4390_/X _4405_/X _4390_/X _4405_/X _4416_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_5396_ _6005_/A _6005_/B _5396_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_160_556 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1011 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1071 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_1150 VGND VPWR sky130_fd_sc_hd__decap_8
X_7135_ _7078_/X _7134_/X _7114_/X _7135_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_4347_ _4345_/X _4346_/X _4344_/X _4347_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_99_684 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_143_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_1149 VGND VPWR sky130_fd_sc_hd__decap_8
X_7066_ _7064_/Y _7065_/Y _7064_/Y _7065_/Y _7066_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_4278_ _4561_/A _4596_/B _4279_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_87_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_902 VGND VPWR sky130_fd_sc_hd__decap_12
X_6017_ _5050_/X _6016_/Y _6017_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_100_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_916 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_426 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_990 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_117 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_269 VGND VPWR sky130_fd_sc_hd__decap_12
X_6919_ _7652_/Q la_data_in[50] _6857_/X _6919_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XPHY_2414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_459 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1001 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1195 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_150 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_684 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_68 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_464 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_68 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_1108 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_183_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_851 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_767 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_846 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_367 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_849 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1207 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_415 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_595 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_286 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_80 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_781 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_932 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1224 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_1115 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1243 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_667 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_121 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_542 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_154_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_872 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_821 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_182_681 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_832 VGND VPWR sky130_fd_sc_hd__decap_12
X_5250_ _5231_/X _5239_/X _5231_/X _5239_/X _5250_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_47_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_142_556 VGND VPWR sky130_fd_sc_hd__decap_12
X_4201_ _4109_/X _4152_/X _4153_/X _4201_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_138_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1233 VGND VPWR sky130_fd_sc_hd__fill_1
X_5181_ _5176_/X _5180_/X _5179_/X _5181_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_190_1252 VGND VPWR sky130_fd_sc_hd__decap_12
X_4132_ _4132_/A _4132_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_3_62 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_1258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_816 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1269 VGND VPWR sky130_fd_sc_hd__decap_8
X_4063_ _4051_/X _4059_/X _4063_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_56_529 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_721 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_497 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_337 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1035 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_384 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_395 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_551 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_916 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_1048 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1056 VGND VPWR sky130_fd_sc_hd__decap_12
X_7753_ _7753_/D _7753_/Q _7797_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_178_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_729 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_459 VGND VPWR sky130_fd_sc_hd__decap_12
X_4965_ _4409_/X _4410_/X _4409_/X _4410_/X _4965_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6704_ _6644_/X _6702_/X _6703_/Y _6704_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XPHY_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_239 VGND VPWR sky130_fd_sc_hd__decap_12
X_3916_ _4959_/A _4583_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_178_954 VGND VPWR sky130_fd_sc_hd__decap_12
X_7684_ _6704_/X _7684_/Q _7707_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4896_ _4479_/B _4898_/D VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_177_453 VGND VPWR sky130_fd_sc_hd__decap_12
X_6635_ _6635_/A _6634_/Y _6635_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_137_306 VGND VPWR sky130_fd_sc_hd__decap_12
X_3847_ _3846_/X _3838_/B _3847_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_20_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_118_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1081 VGND VPWR sky130_fd_sc_hd__decap_12
X_6566_ _6550_/X _6565_/X _6481_/X _6566_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_3778_ _3778_/A _4513_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_180_607 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1062 VGND VPWR sky130_fd_sc_hd__decap_12
X_5517_ _5516_/X _5518_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_106_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_501 VGND VPWR sky130_fd_sc_hd__decap_12
X_6497_ _6495_/Y _6496_/Y _6497_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_5448_ _5383_/Y _5384_/X _5383_/Y _5384_/X _5448_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_195_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1158 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_729 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_910 VGND VPWR sky130_fd_sc_hd__decap_12
X_5379_ _5337_/X _5358_/X _5337_/X _5358_/X _5379_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_120_239 VGND VPWR sky130_fd_sc_hd__decap_12
X_7118_ _7128_/A _7118_/B _7117_/Y _7118_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_59_367 VGND VPWR sky130_fd_sc_hd__decap_12
X_7049_ _7627_/Q _7049_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_74_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1074 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_754 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_819 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_702 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1254 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_70_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_757 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_163_1129 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_151_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_932 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_571 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_328 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_531 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1124 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_372 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1203 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_832 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1236 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_556 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_375 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_698 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_849 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1250 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_326 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_743 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_1125 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1015 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_209_1026 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_1248 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_179_729 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_1207 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_245 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_178_239 VGND VPWR sky130_fd_sc_hd__decap_12
X_4750_ _4748_/X _4749_/X _4750_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_3490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_930 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1013 VGND VPWR sky130_fd_sc_hd__decap_4
X_3701_ wbs_adr_i[16] wbs_adr_i[19] wbs_adr_i[18] wbs_adr_i[21] _3707_/A VGND VPWR
+ sky130_fd_sc_hd__or4_4
XFILLER_159_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_913 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_202_571 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_306 VGND VPWR sky130_fd_sc_hd__decap_8
X_4681_ _4679_/X _4680_/X _4681_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_6420_ _6418_/Y _6420_/B _6420_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_174_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_1158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_618 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_350 VGND VPWR sky130_fd_sc_hd__decap_12
X_6351_ _6333_/A _6354_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_190_938 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_115_501 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_383 VGND VPWR sky130_fd_sc_hd__decap_12
X_5302_ _5300_/X _5301_/X _5532_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_115_534 VGND VPWR sky130_fd_sc_hd__decap_12
X_6282_ _6240_/A _6282_/B _6281_/X _6282_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_89_919 VGND VPWR sky130_fd_sc_hd__decap_12
X_5233_ _5233_/A _4455_/B _5233_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_9_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_1172 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_190_1060 VGND VPWR sky130_fd_sc_hd__decap_8
X_5164_ _5162_/X _5163_/X _5164_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_116_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_1036 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_762 VGND VPWR sky130_fd_sc_hd__decap_12
X_4115_ _4844_/A _4499_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_96_473 VGND VPWR sky130_fd_sc_hd__decap_12
X_5095_ _5095_/A _4903_/B _5096_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_99_1137 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_1099 VGND VPWR sky130_fd_sc_hd__decap_8
X_4046_ _3738_/X _4078_/B _4046_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_17_38 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_702 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_532 VGND VPWR sky130_fd_sc_hd__decap_12
X_7805_ _3816_/Y _7805_/Q _7806_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_207 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_526 VGND VPWR sky130_fd_sc_hd__decap_12
X_5997_ _5993_/C _5996_/Y _5997_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XPHY_229 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_15 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_1001 VGND VPWR sky130_fd_sc_hd__fill_1
X_7736_ _7736_/D _4289_/A _7801_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_40_738 VGND VPWR sky130_fd_sc_hd__decap_12
X_4948_ _7773_/Q _4949_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_149_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_48 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1151 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_952 VGND VPWR sky130_fd_sc_hd__decap_12
X_7667_ _6815_/X _6748_/A _7658_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_166_935 VGND VPWR sky130_fd_sc_hd__decap_8
X_4879_ _4877_/X _4878_/X _4877_/X _4878_/X _4879_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_149_59 VGND VPWR sky130_fd_sc_hd__fill_2
X_6618_ _7690_/Q _6618_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_7598_ _7598_/HI la_data_out[125] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_137_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1269 VGND VPWR sky130_fd_sc_hd__decap_8
X_6549_ _6504_/Y _6505_/Y _6506_/X _6548_/X _6549_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_118_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_639 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_116 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_180_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_898 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_930 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1242 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_67 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_762 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_199_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_359 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_551 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_638 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_128_1002 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_245 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_373 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_203_379 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_913 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_440 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_581 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_141_1235 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_637 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_934 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_434 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_810 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_171_426 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_320 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1085 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_504 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_922 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_996 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_304 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1110 VGND VPWR sky130_fd_sc_hd__decap_8
X_5920_ _7750_/Q _5920_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_0_63 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_841 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_532 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_207_696 VGND VPWR sky130_fd_sc_hd__decap_12
X_5851_ _5841_/X _5842_/X _5841_/X _5842_/X _5851_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_179_515 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_1018 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_727 VGND VPWR sky130_fd_sc_hd__decap_12
X_4802_ _4737_/X _4791_/X _4800_/X _4801_/X _4802_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_5782_ _5757_/X _5758_/X _5757_/X _5758_/X _5782_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_61_395 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_203_880 VGND VPWR sky130_fd_sc_hd__decap_8
X_7521_ _7521_/HI la_data_out[48] VGND VPWR sky130_fd_sc_hd__conb_1
X_4733_ _4712_/X _4730_/X _4731_/X _4732_/X _4733_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_148_935 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_760 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_83 VGND VPWR sky130_fd_sc_hd__decap_8
X_7452_ _7452_/HI io_out[17] VGND VPWR sky130_fd_sc_hd__conb_1
X_4664_ _4664_/A _4665_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_119_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_776 VGND VPWR sky130_fd_sc_hd__decap_12
X_6403_ _7721_/Q _6403_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_147_489 VGND VPWR sky130_fd_sc_hd__decap_12
X_7383_ io_in[30] _7383_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_134_117 VGND VPWR sky130_fd_sc_hd__decap_12
X_4595_ _4512_/A _4595_/B _4595_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_116_832 VGND VPWR sky130_fd_sc_hd__decap_12
X_6334_ _4078_/B _6334_/B _6336_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_162_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_813 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_898 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108 VGND VPWR sky130_fd_sc_hd__decap_12
X_6265_ _6265_/A _6264_/X _7759_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_88_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_548 VGND VPWR sky130_fd_sc_hd__fill_1
X_5216_ _5216_/A _3938_/A _5216_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_6196_ _6089_/X _6193_/X _6195_/X _7770_/D VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_9_1074 VGND VPWR sky130_fd_sc_hd__fill_1
X_5147_ _5146_/A _5146_/B _5146_/X _5147_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_111_570 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_410 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_326 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_151_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_123 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_454 VGND VPWR sky130_fd_sc_hd__decap_4
X_5078_ _4665_/A _4847_/B _5078_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_56_178 VGND VPWR sky130_fd_sc_hd__decap_6
X_4029_ _7784_/Q _4029_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_53_852 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_924 VGND VPWR sky130_fd_sc_hd__fill_2
X_7719_ _7719_/D _6409_/A _7785_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_178_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_1118 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_1011 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_776 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_193_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_467 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_154_938 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_162_971 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_662 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_708 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_664 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_613 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_928 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_958 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_841 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_633 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_874 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_677 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_1013 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1032 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1057 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_765 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_905 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_145_916 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_89_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_757 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_171_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_459 VGND VPWR sky130_fd_sc_hd__decap_12
X_4380_ _4324_/X _4375_/X _4324_/X _4375_/X _4380_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_125_695 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_334 VGND VPWR sky130_fd_sc_hd__fill_2
X_6050_ _6332_/A _6050_/B _6049_/X _6050_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_140_654 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1011 VGND VPWR sky130_fd_sc_hd__decap_12
X_5001_ _4994_/X _4995_/X _4994_/X _4995_/X _5001_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_66_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1123 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_635 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_1186 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_1145 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1028 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_443 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_1039 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_329 VGND VPWR sky130_fd_sc_hd__decap_6
X_6952_ _6952_/A _6952_/B _6952_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_187_1257 VGND VPWR sky130_fd_sc_hd__decap_12
X_5903_ _5901_/X _5902_/X _5901_/X _5902_/X _5903_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_35_863 VGND VPWR sky130_fd_sc_hd__fill_1
X_6883_ la_data_in[63] _6884_/B _6883_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_50_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_502 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_373 VGND VPWR sky130_fd_sc_hd__decap_12
X_5834_ _5831_/X _5832_/X _5833_/X _5834_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_201_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_844 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_710 VGND VPWR sky130_fd_sc_hd__decap_12
X_5765_ _5765_/A _5765_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_22_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_194_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_743 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1252 VGND VPWR sky130_fd_sc_hd__decap_12
X_4716_ _4716_/A _4665_/B _4716_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7504_ _7504_/HI la_data_out[31] VGND VPWR sky130_fd_sc_hd__conb_1
X_5696_ _5594_/X _5595_/X _5594_/X _5595_/X _5696_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_120_1116 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_590 VGND VPWR sky130_fd_sc_hd__decap_12
X_7435_ io_oeb[30] _7435_/LO VGND VPWR sky130_fd_sc_hd__conb_1
X_4647_ _5162_/A _4647_/B _4647_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_30_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_532 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_194_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_7366_ _5062_/Y _7355_/X _7365_/X wbs_dat_o[18] VGND VPWR sky130_fd_sc_hd__o21ai_4
X_4578_ _4560_/X _4576_/X _4560_/X _4576_/X _4578_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6317_ _3904_/X _5275_/X _6317_/C _6317_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_157_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_513 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_524 VGND VPWR sky130_fd_sc_hd__decap_12
X_7297_ _5894_/A _7280_/X _7292_/X _7296_/Y wbs_dat_o[5] VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_116_695 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_118_1045 VGND VPWR sky130_fd_sc_hd__decap_8
X_6248_ _5993_/D _6247_/X _5996_/Y _6248_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_162_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_1242 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_922 VGND VPWR sky130_fd_sc_hd__decap_12
X_6179_ _4983_/X _6178_/X _6179_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_44_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_808 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_999 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_318 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_690 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_164_1032 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_1095 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_186_849 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_539 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_1062 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_426 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_154_746 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_908 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_662 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_684 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_930 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1044 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_288 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1036 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_703 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_483 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_736 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_616 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_104 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_733 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_424 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_1133 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_852 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_863 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_479 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_885 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_182_1121 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_964 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1203 VGND VPWR sky130_fd_sc_hd__decap_12
X_3880_ _3757_/A _3897_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_43_192 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_177_838 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_337 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_390 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_220 VGND VPWR sky130_fd_sc_hd__decap_12
X_5550_ _5543_/X _5544_/X _5543_/X _5544_/X _5550_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_118_905 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_157_562 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_318 VGND VPWR sky130_fd_sc_hd__decap_12
X_4501_ _4500_/A _4500_/B _4500_/X _4501_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_117_415 VGND VPWR sky130_fd_sc_hd__decap_12
X_5481_ _4741_/A _4293_/X _5483_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_172_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_297 VGND VPWR sky130_fd_sc_hd__decap_8
X_7220_ _7199_/X _7218_/X _7219_/Y _7220_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA_0 _4459_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_4432_ _4389_/X _4417_/X _4389_/X _4417_/X _4432_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_126_971 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_587 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_99_822 VGND VPWR sky130_fd_sc_hd__decap_12
X_7151_ _7151_/A _7151_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4363_ _4363_/A _4612_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_99_855 VGND VPWR sky130_fd_sc_hd__decap_12
X_6102_ _4108_/B _6099_/X _6101_/X _6102_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_141_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_440 VGND VPWR sky130_fd_sc_hd__decap_3
X_7082_ _7064_/Y _7065_/Y _7130_/B _7083_/B VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_99_888 VGND VPWR sky130_fd_sc_hd__decap_12
X_4294_ _4898_/A _4293_/X _4301_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_141_996 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_304 VGND VPWR sky130_fd_sc_hd__decap_12
X_6033_ _6033_/A _6060_/B _6034_/C VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_98_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_538 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_140_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_730 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_1044 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_763 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1021 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_947 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_755 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_457 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_16 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6935_ _7645_/Q _6935_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_38 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_660 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_27 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_49 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_693 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_912 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_844 VGND VPWR sky130_fd_sc_hd__decap_8
X_6866_ _6866_/A _6865_/X _6866_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_195_602 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_855 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5817_ _5782_/X _5814_/X _5815_/X _5816_/X _5817_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XPHY_1928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_635 VGND VPWR sky130_fd_sc_hd__decap_12
X_6797_ _6760_/X _6796_/X _6785_/X _6797_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XPHY_1939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1249 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_1090 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_398 VGND VPWR sky130_fd_sc_hd__decap_12
X_5748_ _5679_/X _5704_/B _5704_/X _5748_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_157_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1060 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_735 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_426 VGND VPWR sky130_fd_sc_hd__decap_12
X_5679_ _5668_/A _5667_/X _5668_/X _5679_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_157_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_159_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_459 VGND VPWR sky130_fd_sc_hd__decap_12
X_7418_ io_oeb[13] _7418_/LO VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_11_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_7349_ _7370_/A _7349_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_104_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1217 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_462 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_700 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_796 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_733 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_649 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1116 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_468 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_4543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_479 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_276 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_129 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_181 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_934 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_354 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_158_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1130 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_713 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_971 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_825 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_996 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_730 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_280 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_522 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_533 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_679 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_1206 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_555 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_413 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_566 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_210 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_1227 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_563 VGND VPWR sky130_fd_sc_hd__decap_12
X_4981_ _4982_/A _4982_/B _6015_/A VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_23_107 VGND VPWR sky130_fd_sc_hd__decap_12
X_3932_ _4217_/B _3950_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_6720_ _6720_/A _6720_/B _6720_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_108_1000 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_205_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_192 VGND VPWR sky130_fd_sc_hd__decap_12
X_6651_ _6624_/Y _6625_/Y _6626_/X _6650_/X _6651_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_3863_ _5072_/A _3838_/B _3865_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_149_326 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_825 VGND VPWR sky130_fd_sc_hd__decap_12
X_5602_ _5602_/A _4493_/X _5602_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_31_184 VGND VPWR sky130_fd_sc_hd__decap_12
X_6582_ _7704_/Q la_data_in[6] _6518_/X _6582_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_192_605 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1252 VGND VPWR sky130_fd_sc_hd__decap_12
X_3794_ _4771_/A _4554_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_176_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_1105 VGND VPWR sky130_fd_sc_hd__decap_12
X_5533_ _3738_/X _5533_/B _5533_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_121_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_380 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_245 VGND VPWR sky130_fd_sc_hd__decap_12
X_5464_ _5416_/X _5417_/X _5418_/X _5464_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_105_418 VGND VPWR sky130_fd_sc_hd__decap_8
X_7203_ _7144_/X _7203_/B _7203_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_172_373 VGND VPWR sky130_fd_sc_hd__decap_12
X_4415_ _4411_/X _4414_/X _4411_/X _4414_/X _4415_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_132_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_5395_ _5286_/X _5287_/X _5286_/X _5287_/X _6005_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_99_630 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1023 VGND VPWR sky130_fd_sc_hd__decap_12
X_7134_ _7070_/A la_data_in[82] _7072_/X _7134_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_160_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_62 VGND VPWR sky130_fd_sc_hd__decap_12
X_4346_ _4494_/A _4346_/B _4346_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_8_1128 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_1067 VGND VPWR sky130_fd_sc_hd__fill_1
X_7065_ la_data_in[84] _7065_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_4277_ _4277_/A _4596_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_143_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_657 VGND VPWR sky130_fd_sc_hd__decap_12
X_6016_ _6012_/Y _6013_/X _6015_/X _6016_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_189_1127 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1234 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_914 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_711 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_703 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_3105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_928 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_3116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_276 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_747 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_438 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_129 VGND VPWR sky130_fd_sc_hd__decap_4
X_6918_ _6864_/X _6916_/X _6917_/Y _6918_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XPHY_2415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1100 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_161_1013 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6849_ _7654_/Q _6849_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_1725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_808 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_335 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_476 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_510 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_202_1065 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_779 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_930 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_760 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_172_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_922 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_292 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_390 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_1219 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_93_98 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_298 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_4373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_900 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1203 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1143 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_410 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_944 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_144_1233 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_1236 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1206 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_977 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1228 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_184 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_182_693 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_1026 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_844 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_177_1097 VGND VPWR sky130_fd_sc_hd__fill_1
X_4200_ _4200_/A _4200_/B _4200_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_142_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1220 VGND VPWR sky130_fd_sc_hd__decap_12
X_5180_ _5177_/X _5178_/X _5179_/X _5180_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_4131_ _4131_/A _4127_/X _4132_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_190_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_1237 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_977 VGND VPWR sky130_fd_sc_hd__decap_12
X_4062_ _4040_/X _4061_/X _4040_/X _4061_/X _4062_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_209_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1021 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_850 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_1002 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_149_1122 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_1054 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_703 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_1182 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_872 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_563 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_405 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_276 VGND VPWR sky130_fd_sc_hd__decap_8
X_4964_ _4923_/X _4927_/X _4926_/X _4964_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_7752_ _7752_/D _5867_/A _7797_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_178_922 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_257 VGND VPWR sky130_fd_sc_hd__fill_2
X_6703_ _6644_/X _6702_/X _6690_/X _6703_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_3915_ _4824_/A _4959_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_189_281 VGND VPWR sky130_fd_sc_hd__decap_12
X_4895_ _4485_/B _4959_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_7683_ _6706_/X _7683_/Q _7658_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_149_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_966 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_903 VGND VPWR sky130_fd_sc_hd__decap_12
X_3846_ _4695_/A _3846_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_6634_ la_data_in[19] _6634_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_177_465 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_999 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_318 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_666 VGND VPWR sky130_fd_sc_hd__decap_12
X_3777_ _7809_/Q _3778_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_6565_ _6498_/A la_data_in[12] _6500_/X _6565_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_118_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1093 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_192_457 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_195_1120 VGND VPWR sky130_fd_sc_hd__decap_8
X_5516_ _5516_/A _5516_/B _5516_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_173_660 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_180_619 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1074 VGND VPWR sky130_fd_sc_hd__decap_12
X_6496_ la_data_in[13] _6496_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_106_727 VGND VPWR sky130_fd_sc_hd__decap_12
X_5447_ _5435_/X _5436_/X _5434_/X _5437_/X _5447_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_161_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_5378_ _5374_/X _5377_/X _5374_/X _5377_/X _5378_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_87_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_922 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_398 VGND VPWR sky130_fd_sc_hd__decap_12
X_4329_ _4771_/A _4647_/B _4331_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_7117_ _7117_/A _7088_/X _7117_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_113_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_335 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_806 VGND VPWR sky130_fd_sc_hd__decap_12
X_7048_ _7048_/A _7048_/B _7048_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_86_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_349 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_167_1200 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_511 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_86 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_900 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_544 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_769 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1252 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_944 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_994 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_611 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_977 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_583 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_154 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_435 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_830 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1245 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_170_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_384 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_844 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_1248 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_292 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_625 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_338 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_733 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_168_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_755 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_522 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_1219 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1060 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_1071 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1041 VGND VPWR sky130_fd_sc_hd__fill_1
X_3700_ _3700_/A _3699_/X _3700_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_109_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_942 VGND VPWR sky130_fd_sc_hd__decap_4
X_4680_ _4680_/A _4657_/B _4680_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_186_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_159_476 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_174_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_841 VGND VPWR sky130_fd_sc_hd__decap_12
X_6350_ _6350_/A _6350_/B _6349_/Y _6350_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_127_362 VGND VPWR sky130_fd_sc_hd__decap_4
X_5301_ _4844_/A _5301_/B _5301_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_6281_ _6280_/A _6279_/Y _6281_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_143_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_546 VGND VPWR sky130_fd_sc_hd__decap_3
X_5232_ _5176_/A _4747_/B _5232_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_170_674 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_398 VGND VPWR sky130_fd_sc_hd__decap_12
X_5163_ _4655_/A _4758_/B _5163_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_9_1245 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_430 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_1195 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_806 VGND VPWR sky130_fd_sc_hd__decap_12
X_4114_ _4498_/A _3950_/B _4114_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_68_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1097 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_774 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_305 VGND VPWR sky130_fd_sc_hd__decap_12
X_5094_ _5130_/A _5129_/B _5096_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_96_485 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_1149 VGND VPWR sky130_fd_sc_hd__decap_8
X_4045_ _4044_/A _4043_/X _4044_/X _4045_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_83_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_714 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_202 VGND VPWR sky130_fd_sc_hd__decap_12
X_7804_ _3823_/Y _7804_/Q _7806_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_393 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_544 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_208 VGND VPWR sky130_fd_sc_hd__decap_3
X_5996_ _5723_/X _5765_/Y _5995_/X _5996_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XPHY_219 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_197_538 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_886 VGND VPWR sky130_fd_sc_hd__decap_12
X_7735_ _7735_/D _4295_/A _7801_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4947_ _4894_/X _4910_/X _4893_/X _4911_/X _4947_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_149_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1163 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_700 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1166 VGND VPWR sky130_fd_sc_hd__decap_12
X_7666_ _7666_/D _7666_/Q _7658_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_32_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_964 VGND VPWR sky130_fd_sc_hd__decap_12
X_4878_ _4691_/X _4709_/X _4587_/X _4710_/X _4878_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_71_1068 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_638 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_733 VGND VPWR sky130_fd_sc_hd__decap_6
X_6617_ _6615_/Y _6616_/Y _6615_/Y _6616_/Y _6617_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_123_1158 VGND VPWR sky130_fd_sc_hd__fill_1
X_3829_ _4665_/A _4747_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_119_841 VGND VPWR sky130_fd_sc_hd__decap_12
X_7597_ _7597_/HI la_data_out[124] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_181_906 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_800 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_874 VGND VPWR sky130_fd_sc_hd__fill_1
X_6548_ _6507_/Y _6508_/Y _6576_/B _6548_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_192_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_811 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_682 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_165_59 VGND VPWR sky130_fd_sc_hd__fill_2
X_6479_ _7717_/Q la_data_in[115] _6417_/X _6479_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_82_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_79 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_1107 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_485 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_210_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_861 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_563 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_393 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_190 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_717 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_599 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_44 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_931 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1252 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_251 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_452 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1247 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_649 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_446 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_232 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_1042 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_1026 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_640 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_1097 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_1048 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_516 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_953 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_934 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_839 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_316 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_541 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1164 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_1006 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_75 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_853 VGND VPWR sky130_fd_sc_hd__decap_12
X_5850_ _5847_/X _5849_/X _5847_/X _5849_/X _5850_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_0_97 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_185_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_886 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_577 VGND VPWR sky130_fd_sc_hd__decap_3
X_4801_ _4737_/X _4791_/X _4737_/X _4791_/X _4801_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_21_205 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_739 VGND VPWR sky130_fd_sc_hd__decap_12
X_5781_ _5760_/X _5761_/X _5760_/X _5761_/X _5781_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7520_ _7520_/HI la_data_out[47] VGND VPWR sky130_fd_sc_hd__conb_1
X_4732_ _4712_/X _4730_/X _4712_/X _4730_/X _4732_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_148_947 VGND VPWR sky130_fd_sc_hd__decap_12
X_4663_ _4653_/X _4659_/X _4653_/X _4659_/X _4663_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7451_ _7451_/HI io_out[16] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_190_703 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_159 VGND VPWR sky130_fd_sc_hd__decap_12
X_6402_ _6400_/Y _6401_/Y _6400_/Y _6401_/Y _6467_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_163_928 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_788 VGND VPWR sky130_fd_sc_hd__decap_4
X_4594_ _4589_/X _4593_/X _4592_/X _4594_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_7382_ _4529_/Y _7354_/X _7381_/X wbs_dat_o[23] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_174_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_1191 VGND VPWR sky130_fd_sc_hd__decap_12
X_6333_ _6333_/A _6350_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_157_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_844 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1205 VGND VPWR sky130_fd_sc_hd__decap_8
X_6264_ _5503_/Y _6091_/X _6208_/A _6264_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_192_1145 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_825 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_143_696 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_227 VGND VPWR sky130_fd_sc_hd__decap_12
X_5215_ _5215_/A _4217_/B _5215_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_192_1189 VGND VPWR sky130_fd_sc_hd__fill_1
X_6195_ _4580_/Y _6158_/X _6194_/X _6195_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_69_441 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_761 VGND VPWR sky130_fd_sc_hd__decap_12
X_5146_ _5146_/A _5146_/B _5146_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_97_794 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_485 VGND VPWR sky130_fd_sc_hd__decap_3
X_5077_ _5072_/X _5076_/X _5075_/X _5077_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_151_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_1170 VGND VPWR sky130_fd_sc_hd__decap_12
X_4028_ _3956_/X _4027_/X _4028_/X VGND VPWR sky130_fd_sc_hd__xor2_4
XFILLER_53_820 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_672 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_201_818 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_385 VGND VPWR sky130_fd_sc_hd__decap_12
X_5979_ _5954_/X _5963_/X _5978_/X _5979_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_12_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_379 VGND VPWR sky130_fd_sc_hd__decap_12
X_7718_ _6478_/X _6412_/A _7785_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_205_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_593 VGND VPWR sky130_fd_sc_hd__decap_12
X_7649_ _7649_/D io_out[4] _7756_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_165_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1034 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_822 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_490 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_983 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_825 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_621 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_912 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_676 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_923 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_625 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_658 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_135 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_157 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_937 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_414 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_1254 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_814 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_853 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_689 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1063 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_197_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_1025 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_180_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_552 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_608 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_1069 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_777 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_939 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_287 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_663 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_471 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_481 VGND VPWR sky130_fd_sc_hd__decap_6
X_5000_ _4996_/X _4999_/X _4996_/X _4999_/X _5000_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_85_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_912 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_1023 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_3 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_1162 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_794 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_809 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_1168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_617 VGND VPWR sky130_fd_sc_hd__decap_12
X_6951_ la_data_in[70] _6952_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_82_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1269 VGND VPWR sky130_fd_sc_hd__decap_8
X_5902_ _5867_/Y _5868_/X _5867_/Y _5868_/X _5902_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_46_190 VGND VPWR sky130_fd_sc_hd__decap_12
X_6882_ io_out[3] _6881_/X _6884_/B VGND VPWR sky130_fd_sc_hd__xnor2_4
XFILLER_50_812 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_886 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_514 VGND VPWR sky130_fd_sc_hd__decap_4
X_5833_ _5831_/X _5832_/X _5833_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_195_806 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_856 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_379 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_195_828 VGND VPWR sky130_fd_sc_hd__decap_12
X_5764_ _5764_/A _5765_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_148_722 VGND VPWR sky130_fd_sc_hd__decap_12
X_7503_ _7503_/HI la_data_out[30] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_194_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_1136 VGND VPWR sky130_fd_sc_hd__decap_8
X_4715_ _4695_/X _4699_/X _4695_/X _4699_/X _4715_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_148_755 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_1264 VGND VPWR sky130_fd_sc_hd__decap_12
X_5695_ _5680_/X _5686_/X _5693_/X _5694_/X _5695_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_120_1128 VGND VPWR sky130_fd_sc_hd__fill_1
X_7434_ io_oeb[29] _7434_/LO VGND VPWR sky130_fd_sc_hd__conb_1
X_4646_ _4646_/A _5162_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_162_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_449 VGND VPWR sky130_fd_sc_hd__decap_8
X_4577_ _4502_/X _4508_/X _4496_/X _4509_/X _4577_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_7365_ _5069_/A _7349_/X _7363_/Y _7364_/X _7365_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_6316_ _7746_/Q _6316_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_144_994 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_131_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_825 VGND VPWR sky130_fd_sc_hd__decap_4
X_7296_ _5072_/A _7293_/X _7295_/X _7296_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_157_1062 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_536 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_15 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_157_1095 VGND VPWR sky130_fd_sc_hd__decap_3
X_6247_ _5724_/X _5766_/X _6247_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_162_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_130_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_934 VGND VPWR sky130_fd_sc_hd__decap_12
X_6178_ _4988_/Y _6177_/X _6178_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_170_1262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_580 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_293 VGND VPWR sky130_fd_sc_hd__decap_12
X_5129_ _4771_/A _5129_/B _5129_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_131_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_263 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_820 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_4714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_330 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_514 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_164_1044 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_604 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_198_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_491 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1252 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1074 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_928 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_265 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_713 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_201 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_758 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_419 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_1083 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_942 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1176 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_1195 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_666 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_495 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_748 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_820 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_1145 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_806 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_699 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_380 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_176_349 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_391 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_809 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_232 VGND VPWR sky130_fd_sc_hd__decap_12
X_4500_ _4500_/A _4500_/B _4500_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_5480_ _3846_/X _4366_/B _5480_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_172_511 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_144_202 VGND VPWR sky130_fd_sc_hd__decap_12
X_4431_ _4420_/X _4430_/X _4420_/X _4430_/X _4431_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_172_544 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_1 _4596_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1221 VGND VPWR sky130_fd_sc_hd__decap_12
X_4362_ _4361_/Y _4363_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_7150_ _7150_/A _7150_/B _7150_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_98_300 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_834 VGND VPWR sky130_fd_sc_hd__decap_12
X_6101_ _6308_/B _6101_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_7081_ _7066_/X _7081_/B _7130_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_99_867 VGND VPWR sky130_fd_sc_hd__fill_2
X_4293_ _4570_/B _4293_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_141_964 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_154 VGND VPWR sky130_fd_sc_hd__decap_12
X_6032_ _3993_/Y _4036_/Y _6031_/Y _6060_/B VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_100_316 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_937 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1033 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_639 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_17 VGND VPWR sky130_fd_sc_hd__decap_3
X_6934_ _6934_/A _6934_/B _6934_/X VGND VPWR sky130_fd_sc_hd__and2_4
XPHY_3309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_28 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_39 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_992 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_2619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1236 VGND VPWR sky130_fd_sc_hd__decap_12
X_6865_ _6852_/Y _6853_/Y _6854_/X _6864_/X _6865_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_211_924 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_50_642 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_867 VGND VPWR sky130_fd_sc_hd__decap_12
X_5816_ _5782_/X _5814_/X _5782_/X _5814_/X _5816_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_1918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6796_ _7673_/Q la_data_in[39] _6732_/X _6796_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_167_338 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_647 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1203 VGND VPWR sky130_fd_sc_hd__decap_12
X_5747_ _5727_/X _5746_/X _5747_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_136_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_928 VGND VPWR sky130_fd_sc_hd__decap_12
X_5678_ _5673_/X _5674_/X _5673_/X _5674_/X _5678_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_136_747 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_438 VGND VPWR sky130_fd_sc_hd__decap_12
X_7417_ io_oeb[12] _7417_/LO VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_159_1135 VGND VPWR sky130_fd_sc_hd__decap_12
X_4629_ _4628_/A _4628_/B _4628_/X _4629_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_117_950 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_566 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_600 VGND VPWR sky130_fd_sc_hd__decap_12
X_7348_ _7348_/A _7259_/A _7348_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_190_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_110 VGND VPWR sky130_fd_sc_hd__decap_12
X_7279_ _5946_/A _7257_/X _7274_/X _7278_/Y wbs_dat_o[2] VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_173_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_666 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_496 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_1081 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_861 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1054 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_712 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_403 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_959 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_907 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_1128 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_694 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_806 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_56 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_207_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1123 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_139_574 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_154_511 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_725 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_126_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1134 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_886 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_964 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_761 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_506 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_742 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_292 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_545 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_1218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_1274 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_1168 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_209_578 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_90 VGND VPWR sky130_fd_sc_hd__fill_2
X_4980_ _4946_/X _4979_/X _4946_/X _4979_/X _4982_/B VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_91_575 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_119 VGND VPWR sky130_fd_sc_hd__decap_3
X_3931_ _4647_/B _4217_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_147_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_642 VGND VPWR sky130_fd_sc_hd__decap_8
X_6650_ _6627_/Y _6628_/Y _6696_/B _6650_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_177_625 VGND VPWR sky130_fd_sc_hd__decap_12
X_3862_ _4741_/A _5072_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_189_496 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_141 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_1067 VGND VPWR sky130_fd_sc_hd__fill_1
X_5601_ _5598_/X _5599_/X _5633_/A _5601_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_20_837 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_177_669 VGND VPWR sky130_fd_sc_hd__fill_2
X_6581_ _6543_/X _6579_/X _6580_/Y _6581_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_3793_ _4640_/A _4771_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_31_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1264 VGND VPWR sky130_fd_sc_hd__decap_12
X_5532_ _5532_/A _5532_/B _5532_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_30_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_392 VGND VPWR sky130_fd_sc_hd__decap_4
X_5463_ _5438_/X _5439_/X _5438_/X _5439_/X _5463_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_117_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_577 VGND VPWR sky130_fd_sc_hd__decap_8
X_7202_ _7145_/Y _7147_/B _7147_/X _7201_/X _7203_/B VGND VPWR sky130_fd_sc_hd__o22a_4
X_4414_ _4412_/X _4413_/X _4412_/X _4413_/X _4414_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_172_385 VGND VPWR sky130_fd_sc_hd__decap_12
X_5394_ _5335_/X _5391_/X _5392_/X _5393_/X _6005_/A VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_132_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_642 VGND VPWR sky130_fd_sc_hd__decap_12
X_7133_ _7079_/X _7131_/X _7132_/Y _7133_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_4345_ _4342_/X _4344_/B _4344_/X _4345_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_28_1035 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1005 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_997 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_154_1065 VGND VPWR sky130_fd_sc_hd__decap_3
X_4276_ _4479_/A _4597_/B _4276_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7064_ _7064_/A _7064_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_141_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_859 VGND VPWR sky130_fd_sc_hd__fill_1
X_6015_ _6015_/A _6014_/Y _6015_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_101_669 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1246 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_926 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_403 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_723 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_907 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_609 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_3106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_288 VGND VPWR sky130_fd_sc_hd__decap_6
X_6917_ _6864_/X _6916_/X _6905_/X _6917_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XPHY_3139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1022 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_759 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_2416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1112 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_165_1172 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1066 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_130 VGND VPWR sky130_fd_sc_hd__decap_12
X_6848_ _6846_/Y _6847_/Y _6846_/Y _6847_/Y _6911_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XPHY_2449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_450 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_168_658 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_242 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_483 VGND VPWR sky130_fd_sc_hd__decap_12
X_6779_ _6768_/X _6778_/X _6690_/X _6779_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XPHY_1759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_1022 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_714 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_544 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_163_341 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_555 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_525 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_942 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_934 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_509 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_745 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_907 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_428 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_92_1122 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_4374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_759 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_912 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_93 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_642 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_199_794 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_743 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_220 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1248 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_686 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_123 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_989 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_196 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_166_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_717 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_791 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_170_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1232 VGND VPWR sky130_fd_sc_hd__decap_12
X_4130_ _4112_/X _4129_/X _4112_/X _4129_/X _4130_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_25_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_794 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_190_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_433 VGND VPWR sky130_fd_sc_hd__decap_8
X_4061_ _4041_/X _4047_/X _4048_/X _4060_/X _4061_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_111_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_550 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_561 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_477 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_342 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_1060 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_881 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_353 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1033 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_862 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_575 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_417 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1156 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_92_895 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_1099 VGND VPWR sky130_fd_sc_hd__decap_12
X_7751_ _6298_/Y _5894_/A _7797_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_197_709 VGND VPWR sky130_fd_sc_hd__decap_12
X_4963_ _4918_/X _4919_/X _4917_/X _4963_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_184_1069 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_940 VGND VPWR sky130_fd_sc_hd__decap_8
X_6702_ _7684_/Q la_data_in[18] _6638_/X _6702_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_3914_ _3914_/A _4824_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_178_934 VGND VPWR sky130_fd_sc_hd__decap_12
X_7682_ _7682_/D _6641_/A _7658_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_32_450 VGND VPWR sky130_fd_sc_hd__decap_8
X_4894_ _4840_/X _4848_/X _4839_/X _4849_/X _4894_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_189_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_483 VGND VPWR sky130_fd_sc_hd__decap_8
X_6633_ _6633_/A _6635_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_178_978 VGND VPWR sky130_fd_sc_hd__decap_6
X_3845_ _4749_/A _4695_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_177_477 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_678 VGND VPWR sky130_fd_sc_hd__decap_12
X_6564_ _6551_/X _6562_/X _6563_/Y _6564_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_121_1020 VGND VPWR sky130_fd_sc_hd__decap_12
X_3776_ _3769_/A _3774_/X _3775_/Y _3776_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_118_544 VGND VPWR sky130_fd_sc_hd__fill_1
X_5515_ _5462_/X _5512_/X _5513_/X _5514_/X _5516_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_145_330 VGND VPWR sky130_fd_sc_hd__fill_1
X_6495_ _6495_/A _6495_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_146_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_1105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_160_300 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_739 VGND VPWR sky130_fd_sc_hd__decap_12
X_5446_ _5442_/X _5444_/X _5507_/A _5445_/Y _5446_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_161_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_709 VGND VPWR sky130_fd_sc_hd__decap_12
X_5377_ _5375_/X _5376_/X _5375_/X _5376_/X _5377_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_59_303 VGND VPWR sky130_fd_sc_hd__fill_2
X_7116_ _7090_/X _7113_/X _7115_/Y _7116_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_87_623 VGND VPWR sky130_fd_sc_hd__decap_3
X_4328_ _5128_/A _4328_/B _4328_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_102_934 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_347 VGND VPWR sky130_fd_sc_hd__decap_12
X_7047_ la_data_in[90] _7048_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_75_818 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1010 VGND VPWR sky130_fd_sc_hd__fill_1
X_4259_ _4220_/X _4221_/X _4220_/X _4221_/X _4259_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_86_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_881 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_531 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1212 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_350 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_394 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_912 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_187_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_556 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_422 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_956 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_540 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_781 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_204_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_623 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_196_764 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_488 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_959 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_691 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_166 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_447 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_842 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_188 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_164_661 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_152_856 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_855 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_794 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_398 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_764 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_678 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_775 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_306 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_1252 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_637 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1274 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_206_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_767 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_501 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_288 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_160_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_179_709 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_534 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_940 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1050 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_18_1001 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_4182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_450 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1083 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_1067 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1048 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_1250 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1234 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_853 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_672 VGND VPWR sky130_fd_sc_hd__decap_12
X_5300_ _4570_/A _5300_/B _5300_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_52_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_6280_ _6280_/A _6279_/Y _6282_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_6_682 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_333 VGND VPWR sky130_fd_sc_hd__decap_3
X_5231_ _5218_/X _5219_/X _5218_/X _5219_/X _5231_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_103_709 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_1202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_686 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_623 VGND VPWR sky130_fd_sc_hd__decap_6
X_5162_ _5162_/A _4757_/B _5162_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_25_1038 VGND VPWR sky130_fd_sc_hd__decap_4
X_4113_ _4077_/X _4078_/X _4077_/X _4078_/X _4113_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_57_818 VGND VPWR sky130_fd_sc_hd__decap_12
X_5093_ _5052_/A _4906_/B _5093_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_116_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_317 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_497 VGND VPWR sky130_fd_sc_hd__decap_12
X_4044_ _4044_/A _4043_/X _4044_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_83_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_726 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_586 VGND VPWR sky130_fd_sc_hd__decap_12
X_7803_ _3832_/Y _3826_/A _7806_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_5995_ _5721_/Y _5722_/Y _5995_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_209 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_169_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_556 VGND VPWR sky130_fd_sc_hd__decap_12
X_7734_ _7734_/D _4361_/A _7801_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4946_ _4885_/X _4889_/X _4891_/X _4946_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_80_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_1194 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_792 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_178_764 VGND VPWR sky130_fd_sc_hd__decap_8
X_7665_ _7665_/D io_out[3] _7758_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4877_ _4817_/X _4876_/X _4817_/X _4876_/X _4877_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_149_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_1175 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_712 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1126 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_1178 VGND VPWR sky130_fd_sc_hd__decap_12
X_6616_ la_data_in[25] _6616_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_165_425 VGND VPWR sky130_fd_sc_hd__fill_2
X_3828_ _4548_/A _4665_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_166_959 VGND VPWR sky130_fd_sc_hd__decap_12
X_7596_ _7596_/HI la_data_out[123] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_20_475 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_203_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_609 VGND VPWR sky130_fd_sc_hd__fill_1
X_6547_ _6575_/A _6546_/X _6576_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_3759_ _3759_/A _3790_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_165_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_146_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_385 VGND VPWR sky130_fd_sc_hd__decap_12
X_6478_ _6466_/X _6429_/X _6477_/Y _6478_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_5429_ _5428_/A _5427_/X _5428_/X _5431_/A VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_160_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_528 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_825 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_1154 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_869 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_1187 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_306 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_1119 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_648 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_1154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_629 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_501 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_575 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_692 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_517 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1097 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_729 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_56 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_550 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_943 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_11_420 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_701 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_1275 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_105 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_464 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1259 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_947 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_609 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_428 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_178_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_940 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_152_631 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_152_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1133 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_174_1024 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_630 VGND VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_1_1_1_wb_clk_i clkbuf_1_1_0_wb_clk_i/X clkbuf_1_1_1_wb_clk_i/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_3_652 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_729 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_1188 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_965 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_818 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_328 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_1121 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_840 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1093 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_0_0_wb_clk_i clkbuf_3_0_0_wb_clk_i/X _7658_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_4_1176 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_361 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1018 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_87 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_545 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_865 VGND VPWR sky130_fd_sc_hd__decap_12
X_4800_ _4796_/X _4799_/X _4796_/X _4799_/X _4800_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_94_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_364 VGND VPWR sky130_fd_sc_hd__fill_2
X_5780_ _5775_/X _5779_/X _5993_/C VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_21_217 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_792 VGND VPWR sky130_fd_sc_hd__fill_1
X_4731_ _4542_/X _4543_/X _4542_/X _4543_/X _4731_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_187_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_403 VGND VPWR sky130_fd_sc_hd__fill_2
X_7450_ _7450_/HI io_out[15] VGND VPWR sky130_fd_sc_hd__conb_1
X_4662_ _4644_/X _4661_/X _4644_/X _4661_/X _4662_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_148_959 VGND VPWR sky130_fd_sc_hd__decap_8
X_6401_ la_data_in[120] _6401_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_7381_ _3693_/X _7370_/X _7380_/Y _7265_/X _7381_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_4593_ _4592_/A _4592_/B _4592_/X _4593_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_174_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_300 VGND VPWR sky130_fd_sc_hd__decap_4
X_6332_ _6332_/A _6332_/B _6331_/Y _7744_/D VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_127_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1097 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_322 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_157_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_490 VGND VPWR sky130_fd_sc_hd__decap_12
X_6263_ _6240_/A _6261_/X _6263_/C _6265_/A VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_171_984 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_729 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_192_1157 VGND VPWR sky130_fd_sc_hd__decap_12
X_5214_ _5198_/X _5202_/X _5198_/X _5202_/X _5214_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_88_239 VGND VPWR sky130_fd_sc_hd__decap_12
X_6194_ _6144_/A _6194_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_69_453 VGND VPWR sky130_fd_sc_hd__decap_12
X_5145_ _4666_/A _4844_/B _5146_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_111_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_773 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_604 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1087 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_594 VGND VPWR sky130_fd_sc_hd__fill_1
X_5076_ _5073_/X _5074_/X _5075_/X _5076_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_42_1182 VGND VPWR sky130_fd_sc_hd__decap_8
X_4027_ _3970_/Y _4027_/B _4027_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_38_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_832 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_198_815 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_1215 VGND VPWR sky130_fd_sc_hd__decap_12
X_5978_ _5954_/X _5978_/B _5978_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_7717_ _7717_/D _7717_/Q _7785_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_12_239 VGND VPWR sky130_fd_sc_hd__decap_12
X_4929_ _4392_/X _4396_/X _4392_/X _4396_/X _4929_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_100_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_701 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_712 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1245 VGND VPWR sky130_fd_sc_hd__decap_12
X_7648_ _7648_/D _7648_/Q _7754_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_193_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_7579_ _7579_/HI la_data_out[106] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_101_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_586 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_928 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_153_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_620 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_995 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_686 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_633 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_902 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_1041 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_935 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_637 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_91_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_607 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_1233 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_169 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_169_1148 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_61 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_426 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_1266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_459 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_556 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_203_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_898 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_589 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1020 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_548 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_403 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_93 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1143 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_745 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_261 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_789 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_172_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_940 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_171_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_804 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_601 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_153_995 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1035 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_152_1174 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_732 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_776 VGND VPWR sky130_fd_sc_hd__fill_2
X_6950_ _6950_/A _6952_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_54_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_207_440 VGND VPWR sky130_fd_sc_hd__decap_12
X_5901_ _5897_/X _5900_/X _5901_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_6881_ _6819_/Y _6820_/Y _6880_/X _6881_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_5832_ _3877_/A _4482_/A _5832_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_210_605 VGND VPWR sky130_fd_sc_hd__decap_12
X_5763_ _5725_/X _5762_/X _5764_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_201_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_868 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_559 VGND VPWR sky130_fd_sc_hd__decap_12
X_7502_ _7502_/HI la_data_out[29] VGND VPWR sky130_fd_sc_hd__conb_1
X_4714_ _4701_/X _4702_/X _4701_/X _4702_/X _4714_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_148_734 VGND VPWR sky130_fd_sc_hd__fill_2
X_5694_ _5680_/X _5686_/X _5680_/X _5686_/X _5694_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_124_1276 VGND VPWR sky130_fd_sc_hd__fill_1
X_7433_ io_oeb[28] _7433_/LO VGND VPWR sky130_fd_sc_hd__conb_1
X_4645_ _4645_/A _4653_/B _4645_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_200_1120 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_748 VGND VPWR sky130_fd_sc_hd__decap_12
X_7364_ _7351_/B _7364_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4576_ _4567_/X _4575_/X _4567_/X _4575_/X _4576_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_6315_ _6106_/X _6313_/X _6314_/X _7747_/D VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_116_675 VGND VPWR sky130_fd_sc_hd__fill_1
X_7295_ _7295_/A _7300_/B _7295_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_131_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_548 VGND VPWR sky130_fd_sc_hd__fill_1
X_6246_ _5775_/X _6246_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_115_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_1069 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_358 VGND VPWR sky130_fd_sc_hd__decap_8
X_6177_ _6174_/Y _6176_/X _6177_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_130_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_1252 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_1214 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_170_1274 VGND VPWR sky130_fd_sc_hd__decap_3
X_5128_ _5128_/A _4512_/B _5128_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_111_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_916 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_131_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_5059_ _5059_/A _5059_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_57_489 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_72_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_180 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_4748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_865 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_4759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_971 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_678 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_627 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_570 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_1248 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_1086 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_715 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_181_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_288 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_725 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_14_1081 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1062 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_910 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_984 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_1095 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_1188 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_1038 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_678 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_441 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_924 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_986 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_997 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_716 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_380 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_776 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_832 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_757 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_1157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_204_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_188_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_143_1129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_1189 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_367 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_370 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_381 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_392 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_570 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_541 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_428 VGND VPWR sky130_fd_sc_hd__decap_12
X_4430_ _4430_/A _4429_/X _4430_/X VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA_2 _4830_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_556 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1233 VGND VPWR sky130_fd_sc_hd__decap_12
X_4361_ _4361_/A _4361_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_160_729 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_1203 VGND VPWR sky130_fd_sc_hd__decap_12
X_6100_ _4108_/B _6099_/X _6100_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_113_623 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_846 VGND VPWR sky130_fd_sc_hd__decap_8
X_7080_ _7067_/Y _7068_/Y _7069_/X _7079_/X _7081_/B VGND VPWR sky130_fd_sc_hd__o22a_4
X_4292_ _4830_/B _4570_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_101_818 VGND VPWR sky130_fd_sc_hd__decap_12
X_6031_ _3994_/A _6031_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_86_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_328 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_551 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_404 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_117 VGND VPWR sky130_fd_sc_hd__decap_8
X_6933_ la_data_in[76] _6934_/B VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_18 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_148_1029 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_459 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_29 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_207_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_1215 VGND VPWR sky130_fd_sc_hd__decap_4
X_6864_ _6857_/A _6857_/B _6857_/X _6863_/X _6864_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XPHY_2609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1248 VGND VPWR sky130_fd_sc_hd__decap_3
X_5815_ _5801_/X _5810_/X _5809_/X _5811_/X _5815_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_34_194 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_306 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_654 VGND VPWR sky130_fd_sc_hd__decap_12
X_6795_ _6795_/A _6762_/X _6795_/C _6795_/X VGND VPWR sky130_fd_sc_hd__and3_4
XPHY_1919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_507 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1081 VGND VPWR sky130_fd_sc_hd__fill_2
X_5746_ _5728_/X _5745_/B _5745_/X _5746_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_195_659 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_884 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_715 VGND VPWR sky130_fd_sc_hd__decap_12
X_5677_ _5643_/X _5676_/X _5643_/X _5676_/X _5677_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_157_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_7416_ io_oeb[11] _7416_/LO VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_68_1008 VGND VPWR sky130_fd_sc_hd__decap_8
X_4628_ _4628_/A _4628_/B _4628_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_194_1016 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_759 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_159_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_962 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_578 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_706 VGND VPWR sky130_fd_sc_hd__decap_8
X_7347_ _5507_/A _7388_/A _7343_/X _7346_/Y wbs_dat_o[14] VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_132_910 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_717 VGND VPWR sky130_fd_sc_hd__decap_8
X_4559_ _4551_/X _4557_/X _4551_/X _4557_/X _4559_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_104_612 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_728 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_739 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_173_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_239 VGND VPWR sky130_fd_sc_hd__decap_12
X_7278_ _5198_/A _7262_/X _7277_/X _7278_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_106_32 VGND VPWR sky130_fd_sc_hd__decap_12
X_6229_ _6189_/A _6227_/X _6228_/Y _6229_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_170_1060 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_231 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_776 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_873 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1115 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_724 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_1099 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_4512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_139 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_684 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_161 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_301 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_4589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_68 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_818 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_643 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_654 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_62 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_3899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_95 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_840 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1146 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_556 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_1130 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_710 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_754 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_595 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_426 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_245 VGND VPWR sky130_fd_sc_hd__decap_12
X_3930_ _3930_/A _4647_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_16_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_172 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_204_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_1062 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_149_306 VGND VPWR sky130_fd_sc_hd__decap_12
X_3861_ _5157_/A _4741_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_32_665 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_637 VGND VPWR sky130_fd_sc_hd__decap_12
X_5600_ _5598_/X _5599_/X _5633_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_6580_ _6543_/X _6579_/X _6572_/X _6580_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_82_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_3792_ _7807_/Q _4640_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_5531_ _5523_/X _5524_/X _5529_/X _5530_/X _5531_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_192_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_715 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_1257 VGND VPWR sky130_fd_sc_hd__decap_12
X_5462_ _5450_/X _5451_/X _5450_/X _5451_/X _5462_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7201_ _7150_/A _7150_/B _7150_/X _7200_/X _7201_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_173_887 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_269 VGND VPWR sky130_fd_sc_hd__decap_12
X_4413_ _4345_/X _4346_/X _4345_/X _4346_/X _4413_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_910 VGND VPWR sky130_fd_sc_hd__fill_2
X_5393_ _5335_/X _5391_/X _5335_/X _5391_/X _5393_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7132_ _7079_/X _7131_/X _7114_/X _7132_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_132_239 VGND VPWR sky130_fd_sc_hd__decap_12
X_4344_ _4342_/X _4344_/B _4344_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_193_1071 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_1108 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_762 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1096 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_1047 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_86 VGND VPWR sky130_fd_sc_hd__decap_12
X_7063_ _7061_/Y _7062_/Y _7061_/Y _7062_/Y _7083_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_115_1017 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1069 VGND VPWR sky130_fd_sc_hd__decap_12
X_4275_ _4145_/A _4597_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_119_1186 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_337 VGND VPWR sky130_fd_sc_hd__decap_12
X_6014_ _4982_/X _4987_/X _6014_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_80_1252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_562 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_1258 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_938 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_757 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_768 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6916_ _7653_/Q la_data_in[51] _6854_/X _6916_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XPHY_2406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1034 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_604 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1124 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_6847_ la_data_in[53] _6847_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_1705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_142 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_27 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_1738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6778_ _7679_/Q la_data_in[45] _6714_/X _6778_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XPHY_1749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_254 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_13_0_wb_clk_i clkbuf_3_6_0_wb_clk_i/X _7806_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_183_607 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_211_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_276 VGND VPWR sky130_fd_sc_hd__decap_12
X_5729_ _5681_/X _5685_/X _5681_/X _5685_/X _5729_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_195_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1034 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_148_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_726 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_184_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1089 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_707 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_353 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_876 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_567 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_684 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_729 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1062 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_781 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_548 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_954 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_816 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_1196 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_1038 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1049 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_871 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_562 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_554 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_459 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_919 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_1252 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_1191 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_4331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_204 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_4353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_941 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_4386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_615 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_654 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_440 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_755 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_201_232 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_135 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_2995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_93 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_158_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_813 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_341 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_729 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_7 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_886 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_114_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1099 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_64_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_879 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_123_751 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_1244 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_315 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_935 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_43 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_337 VGND VPWR sky130_fd_sc_hd__decap_12
X_4060_ _4059_/A _4059_/B _4059_/X _4060_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_96_668 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_456 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_87 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_871 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_1001 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_190_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_510 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_1196 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_1027 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_209_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_1038 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_532 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_757 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_727 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_289 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_429 VGND VPWR sky130_fd_sc_hd__decap_12
X_4962_ _4954_/X _4961_/X _4954_/X _4961_/X _4962_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7750_ _7750_/D _7750_/Q _7797_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_3913_ _7310_/A _3913_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_6701_ _6645_/X _6699_/X _6700_/Y _7685_/D VGND VPWR sky130_fd_sc_hd__o21a_4
X_7681_ _6775_/Y io_out[2] _7758_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4893_ _4833_/X _4834_/X _4826_/X _4835_/X _4893_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_20_602 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_771 VGND VPWR sky130_fd_sc_hd__decap_8
X_6632_ _6630_/Y _6631_/Y _6630_/Y _6631_/Y _6647_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_3844_ _4667_/A _4749_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_149_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_916 VGND VPWR sky130_fd_sc_hd__decap_12
X_6563_ _6551_/X _6562_/X _6481_/X _6563_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_158_670 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_177_489 VGND VPWR sky130_fd_sc_hd__decap_12
X_3775_ wbs_dat_i[16] _3790_/B _3775_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_164_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_1032 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_1081 VGND VPWR sky130_fd_sc_hd__decap_12
X_5514_ _5462_/X _5512_/X _5462_/X _5512_/X _5514_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_192_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1114 VGND VPWR sky130_fd_sc_hd__fill_1
X_6494_ _6492_/Y _6493_/Y _6492_/Y _6493_/Y _6560_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_8_190 VGND VPWR sky130_fd_sc_hd__decap_8
X_5445_ _5442_/X _5444_/X _5442_/X _5444_/X _5445_/Y VGND VPWR sky130_fd_sc_hd__a2bb2oi_4
XFILLER_146_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_1158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_145_386 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_191_1019 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_740 VGND VPWR sky130_fd_sc_hd__fill_2
X_5376_ _5265_/X _5266_/X _5265_/X _5266_/X _5376_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_161_879 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_440 VGND VPWR sky130_fd_sc_hd__decap_12
X_7115_ _7090_/X _7113_/X _7114_/X _7115_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_4327_ _4260_/X _4265_/X _4260_/X _4265_/X _4327_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_160_389 VGND VPWR sky130_fd_sc_hd__decap_8
X_7046_ _7628_/Q _7048_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_101_445 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_359 VGND VPWR sky130_fd_sc_hd__decap_6
X_4258_ _4223_/X _4231_/X _4223_/X _4231_/X _4258_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_86_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_489 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_1093 VGND VPWR sky130_fd_sc_hd__decap_12
X_4189_ _4189_/A _4137_/X _4189_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_55_543 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_1099 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_919 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_3_1_wb_clk_i clkbuf_2_3_0_wb_clk_i/X clkbuf_3_7_0_wb_clk_i/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_82_362 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_1210 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_941 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_924 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_1243 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_440 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_59 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_220 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_968 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_211_552 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_635 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_776 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_415 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_184_938 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_668 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1241 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_971 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_673 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_164_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_868 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_345 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_151_367 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_613 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_1061 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_787 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_1242 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_1250 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_990 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_649 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_690 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_852 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_779 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_727 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_204 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_546 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_4172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_952 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_721 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_985 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_3482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_552 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_1095 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_175_905 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_2770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_916 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_495 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_147_629 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_1038 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1246 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_865 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_898 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_155_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_694 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_160 VGND VPWR sky130_fd_sc_hd__decap_6
X_5230_ _5221_/X _5222_/X _5221_/X _5222_/X _5230_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_170_654 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_900 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_518 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_1214 VGND VPWR sky130_fd_sc_hd__decap_6
X_5161_ _4645_/A _4756_/B _5161_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_170_698 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_1172 VGND VPWR sky130_fd_sc_hd__decap_12
X_4112_ _4080_/X _4087_/X _4080_/X _4087_/X _4112_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_97_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_668 VGND VPWR sky130_fd_sc_hd__decap_3
X_5092_ _5066_/X _5067_/X _5066_/X _5067_/X _5092_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_84_605 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_116_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_178 VGND VPWR sky130_fd_sc_hd__decap_12
X_4043_ _5069_/A _3949_/B _4043_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_84_638 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_329 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_209_140 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_554 VGND VPWR sky130_fd_sc_hd__fill_1
X_7802_ _7802_/D _7802_/Q _7806_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_92_682 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_5994_ _5774_/X _5778_/X _5998_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_52_568 VGND VPWR sky130_fd_sc_hd__decap_12
X_4945_ _4941_/X _4942_/X _4943_/X _4944_/X _4982_/A VGND VPWR sky130_fd_sc_hd__o22a_4
X_7733_ _7733_/D _4480_/A _7801_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_178_743 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_220 VGND VPWR sky130_fd_sc_hd__decap_12
X_4876_ _4874_/X _4875_/X _4874_/X _4875_/X _4876_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7664_ _6887_/X _6819_/A _7754_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_162_1187 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_123_1138 VGND VPWR sky130_fd_sc_hd__decap_12
X_3827_ _4453_/A _4548_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_6615_ _6615_/A _6615_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_193_724 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_977 VGND VPWR sky130_fd_sc_hd__decap_12
X_7595_ _7595_/HI la_data_out[122] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_159_990 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_746 VGND VPWR sky130_fd_sc_hd__decap_12
X_6546_ _6510_/Y _6511_/Y _6545_/X _6546_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_20_498 VGND VPWR sky130_fd_sc_hd__decap_3
X_3758_ _5069_/A _3767_/B _3761_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_203_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_971 VGND VPWR sky130_fd_sc_hd__decap_12
X_6477_ _6429_/A _6429_/B _6477_/Y VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_165_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_835 VGND VPWR sky130_fd_sc_hd__decap_12
X_3689_ _3689_/A _4820_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_106_548 VGND VPWR sky130_fd_sc_hd__decap_12
X_5428_ _5428_/A _5427_/X _5428_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_133_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_5359_ _5253_/X _5257_/X _5253_/X _5257_/X _5359_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_581 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_181_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_605 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_102_776 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_476 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_114_32 VGND VPWR sky130_fd_sc_hd__decap_12
X_7029_ _6970_/X _7027_/X _7028_/Y _7029_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_28_532 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_210_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1010 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_727 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_598 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_167_1065 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_855 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_218 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_398 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_141_1205 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_281 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_403 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_735 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_128_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_999 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_476 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_959 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_183_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_768 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_156_459 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1172 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_654 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_805 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_130 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_664 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_174_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_581 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_413 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_11 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_852 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_1188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_1199 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_1026 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_833 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_598 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_206_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_332 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_1168 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_557 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_877 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_159_220 VGND VPWR sky130_fd_sc_hd__decap_12
X_4730_ _4713_/X _4727_/X _4728_/X _4729_/X _4730_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XPHY_3290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_562 VGND VPWR sky130_fd_sc_hd__decap_12
X_4661_ _4652_/X _4660_/X _4652_/X _4660_/X _4661_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_30_785 VGND VPWR sky130_fd_sc_hd__decap_12
X_6400_ _6400_/A _6400_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_7380_ io_in[29] _7380_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_70_1081 VGND VPWR sky130_fd_sc_hd__decap_8
X_4592_ _4592_/A _4592_/B _4592_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_190_716 VGND VPWR sky130_fd_sc_hd__decap_12
X_6331_ wbs_dat_i[14] _6338_/B _6331_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_128_684 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_183_790 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_857 VGND VPWR sky130_fd_sc_hd__decap_12
X_6262_ _5724_/X _6260_/Y _6263_/C VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_157_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_1128 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_170_451 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_996 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_304 VGND VPWR sky130_fd_sc_hd__decap_12
X_5213_ _5204_/X _5205_/X _5204_/X _5205_/X _5213_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_170_484 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_1169 VGND VPWR sky130_fd_sc_hd__decap_12
X_6193_ _4807_/X _6149_/B _6150_/B _6193_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_130_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_741 VGND VPWR sky130_fd_sc_hd__fill_1
X_5144_ _4655_/A _4915_/B _5146_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_96_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_465 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_562 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_785 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_627 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_318 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_947 VGND VPWR sky130_fd_sc_hd__decap_8
X_5075_ _5073_/X _5074_/X _5075_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_85_958 VGND VPWR sky130_fd_sc_hd__decap_12
X_4026_ _3998_/X _4025_/X _4026_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_53_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1227 VGND VPWR sky130_fd_sc_hd__decap_12
X_5977_ _5975_/X _5977_/B _5978_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7716_ _6486_/X _7716_/Q _7785_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_398 VGND VPWR sky130_fd_sc_hd__decap_12
X_4928_ _4923_/X _4927_/X _4923_/X _4927_/X _4928_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_178_551 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_916 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_724 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1257 VGND VPWR sky130_fd_sc_hd__decap_12
X_7647_ _6997_/X _7647_/Q _7754_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4859_ _4852_/X _4858_/X _4852_/X _4858_/X _4859_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_193_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_1003 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_176_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_459 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_165_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_640 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1252 VGND VPWR sky130_fd_sc_hd__decap_6
X_7578_ _7578_/HI la_data_out[105] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_147_971 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_1274 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_598 VGND VPWR sky130_fd_sc_hd__decap_12
X_6529_ la_data_in[2] _6530_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_106_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_440 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_654 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_107_879 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_816 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_1050 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_645 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_197_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1053 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_413 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_689 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_800 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_73 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_991 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_513 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_693 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_449 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_505 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_188_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_376 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_1032 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_702 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_1160 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_251 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_273 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_1188 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_106_1199 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_156_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_172_727 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_176_1109 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_632 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_93 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_166_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_451 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_816 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_516 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1172 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_152_1142 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_79_785 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_1047 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_1058 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_152_1186 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_744 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_958 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_1205 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_931 VGND VPWR sky130_fd_sc_hd__decap_12
X_5900_ _5898_/X _5899_/X _5900_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_207_452 VGND VPWR sky130_fd_sc_hd__decap_12
X_6880_ _6821_/X _6880_/B _6880_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_35_855 VGND VPWR sky130_fd_sc_hd__decap_8
X_5831_ _3867_/Y _4477_/A _5831_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_50_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_398 VGND VPWR sky130_fd_sc_hd__decap_12
X_5762_ _5726_/X _5759_/X _5760_/X _5761_/X _5762_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_210_617 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_1154 VGND VPWR sky130_fd_sc_hd__decap_12
X_7501_ _7501_/HI la_data_out[28] VGND VPWR sky130_fd_sc_hd__conb_1
X_4713_ _4704_/X _4705_/X _4704_/X _4705_/X _4713_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_5693_ _5690_/X _5691_/X _5692_/X _5693_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_202_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_245 VGND VPWR sky130_fd_sc_hd__decap_12
X_4644_ _4639_/X _4643_/X _4639_/X _4643_/X _4644_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7432_ io_oeb[27] _7432_/LO VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_163_705 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_919 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_4575_ _4573_/X _4574_/X _4573_/X _4574_/X _4575_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7363_ io_in[24] _7363_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_200_1154 VGND VPWR sky130_fd_sc_hd__decap_12
X_6314_ _5957_/Y _6256_/B _3743_/A _6314_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_143_440 VGND VPWR sky130_fd_sc_hd__decap_4
X_7294_ io_in[11] _7295_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_143_451 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_1015 VGND VPWR sky130_fd_sc_hd__decap_8
X_6245_ _6219_/X _6243_/X _6244_/X _7762_/D VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_104_849 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_635 VGND VPWR sky130_fd_sc_hd__decap_6
X_6176_ _6013_/X _6176_/B _6176_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_130_178 VGND VPWR sky130_fd_sc_hd__decap_12
X_5127_ _5122_/X _5126_/X _5122_/X _5126_/X _5127_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_85_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_424 VGND VPWR sky130_fd_sc_hd__decap_3
X_5058_ _5058_/A _5533_/B _5058_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_55_27 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_211_1272 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_276 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4009_ _4007_/X _4008_/X _4009_/X VGND VPWR sky130_fd_sc_hd__or2_4
XPHY_4727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_1002 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_877 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_1027 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_197_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_1276 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_187_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_139_757 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_181_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_1093 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_952 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_1003 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_996 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_910 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_175_1175 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_281 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_161_292 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_453 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_871 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_475 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_728 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_497 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_392 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_227 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_1080 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1170 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_844 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_321 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_855 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_204_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_1097 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1233 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_825 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_184 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_398 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_108_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_360 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_188_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_510 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_371 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_185_830 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_379 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_382 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_393 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_553 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_1182 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_3 _4293_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_172_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_963 VGND VPWR sky130_fd_sc_hd__fill_1
X_4360_ _4359_/A _4358_/X _4359_/X _4360_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_113_602 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_996 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_410 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_324 VGND VPWR sky130_fd_sc_hd__decap_12
X_4291_ _4291_/A _4830_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_6030_ _7321_/A _3966_/B _6033_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_113_668 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1070 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_446 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_563 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_703 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_468 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_276 VGND VPWR sky130_fd_sc_hd__decap_12
X_6932_ _6932_/A _6934_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_208_772 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_181 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_19 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_293 VGND VPWR sky130_fd_sc_hd__decap_12
X_6863_ _6858_/Y _6859_/Y _6862_/X _6863_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_179_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_471 VGND VPWR sky130_fd_sc_hd__decap_12
X_5814_ _5803_/X _5804_/X _5812_/X _5813_/X _5814_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_161_1208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_184 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_210_414 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_335 VGND VPWR sky130_fd_sc_hd__fill_1
X_6794_ _6794_/A _6761_/X _6795_/C VGND VPWR sky130_fd_sc_hd__nand2_4
XFILLER_22_346 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_666 VGND VPWR sky130_fd_sc_hd__decap_12
X_5745_ _5728_/X _5745_/B _5745_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_148_532 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1227 VGND VPWR sky130_fd_sc_hd__decap_12
X_5676_ _5664_/X _5675_/X _5664_/X _5675_/X _5676_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_198_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_727 VGND VPWR sky130_fd_sc_hd__fill_1
X_7415_ io_oeb[10] _7415_/LO VGND VPWR sky130_fd_sc_hd__conb_1
X_4627_ _5095_/A _4641_/B _4628_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_191_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_708 VGND VPWR sky130_fd_sc_hd__decap_12
X_4558_ _4459_/X _4463_/X _4462_/X _4558_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_7346_ _4459_/A _7322_/X _7345_/X _7346_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_117_974 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_922 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_996 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_190_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_624 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_9 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_173_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_495 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_1209 VGND VPWR sky130_fd_sc_hd__decap_8
X_4489_ _4488_/Y _5835_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_7277_ _7275_/Y _7300_/B _7277_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_103_123 VGND VPWR sky130_fd_sc_hd__decap_12
X_6228_ _6228_/A _6228_/B _6228_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_44_1020 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_487 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_6159_ _4376_/Y _6158_/X _6144_/X _6159_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_85_541 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_755 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_254 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_788 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_574 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_1127 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_1078 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_32 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_747 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_205_208 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_410 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_825 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_81_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_173 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_184 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_666 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1160 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_85 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_852 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_185_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1035 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_182_800 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_194_660 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_501 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_1158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_568 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_440 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_142_719 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_900 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_410 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_806 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_880 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_722 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_638 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_766 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_928 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_405 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_438 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_1249 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_205_720 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_419 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_931 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_696 VGND VPWR sky130_fd_sc_hd__decap_12
X_3860_ _4697_/A _5157_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_204_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_318 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_147_1096 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_677 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_649 VGND VPWR sky130_fd_sc_hd__decap_12
X_3791_ _3791_/A _3791_/B _3790_/Y _3791_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_188_80 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_190 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_1252 VGND VPWR sky130_fd_sc_hd__decap_12
X_5530_ _5523_/X _5524_/X _5523_/X _5524_/X _5530_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_185_660 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_727 VGND VPWR sky130_fd_sc_hd__decap_12
X_5461_ _5453_/X _5454_/X _5453_/X _5454_/X _5516_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_121_1269 VGND VPWR sky130_fd_sc_hd__decap_8
X_4412_ _4401_/X _4402_/X _4400_/X _4412_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_7200_ _7151_/Y _7152_/Y _7153_/X _7199_/X _7200_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_133_708 VGND VPWR sky130_fd_sc_hd__fill_1
X_5392_ _5386_/X _5387_/X _5385_/X _5388_/X _5392_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_126_760 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_771 VGND VPWR sky130_fd_sc_hd__decap_8
X_4343_ _4612_/A _4460_/B _4344_/B VGND VPWR sky130_fd_sc_hd__or2_4
X_7131_ _7621_/Q la_data_in[83] _7069_/X _7131_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_193_1050 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_281 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_193_1083 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_666 VGND VPWR sky130_fd_sc_hd__decap_4
X_7062_ la_data_in[85] _7062_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_154_1045 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_154 VGND VPWR sky130_fd_sc_hd__decap_12
X_4274_ _4259_/X _4266_/X _4272_/X _4273_/X _4274_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_141_774 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_1059 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_207_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_1198 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_1029 VGND VPWR sky130_fd_sc_hd__decap_8
X_6013_ _4881_/Y _4883_/B _4806_/Y _4883_/X _6013_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_101_649 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_189_1119 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_80_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_254 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_574 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_544 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_591 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_1111 VGND VPWR sky130_fd_sc_hd__decap_8
X_6915_ _6923_/A _6866_/X _6914_/Y _7654_/D VGND VPWR sky130_fd_sc_hd__and3_4
XPHY_3119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_791 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_931 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_2418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_1046 VGND VPWR sky130_fd_sc_hd__decap_12
X_6846_ _6846_/A _6846_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_168_616 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_806 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_1717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_211_745 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_1158 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_154 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_828 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_149_830 VGND VPWR sky130_fd_sc_hd__decap_12
X_6777_ _6694_/X _6770_/X _6776_/Y _7680_/D VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_23_699 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_176 VGND VPWR sky130_fd_sc_hd__decap_8
X_3989_ _3984_/X _3987_/X _3984_/X _3987_/X _3989_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_167_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_349 VGND VPWR sky130_fd_sc_hd__decap_12
X_5728_ _5693_/X _5694_/X _5693_/X _5694_/X _5728_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_210_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_885 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_309 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_148_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_1057 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_5659_ _5465_/X _5477_/X _5478_/X _5659_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_184_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_579 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_163_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_151_505 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_1074 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_110 VGND VPWR sky130_fd_sc_hd__decap_12
X_7329_ _7329_/A _7324_/B _7329_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_137_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_752 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_966 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_977 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_928 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_883 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_894 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_133_86 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_257 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_4332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_60_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_1233 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_4376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_144_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_251 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_666 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_452 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_103 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_446 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_139_351 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_861 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_177_1012 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_155_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_843 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_888 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_516 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_353 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_898 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_181_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_154_398 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_1215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_763 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_903 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_11 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_174_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_327 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_947 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_55 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_349 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_95_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_541 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_1006 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_188_1130 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_769 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_149_1136 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_886 VGND VPWR sky130_fd_sc_hd__fill_2
X_4961_ _4955_/X _4960_/X _4955_/X _4960_/X _4961_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_52_739 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_550 VGND VPWR sky130_fd_sc_hd__decap_12
X_6700_ _6645_/X _6699_/X _6690_/X _6700_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_3912_ _7315_/A _3993_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_32_430 VGND VPWR sky130_fd_sc_hd__fill_1
X_7680_ _7680_/D _6709_/A _7658_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4892_ _4891_/A _4891_/B _4891_/X _4892_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_71_1219 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_975 VGND VPWR sky130_fd_sc_hd__fill_1
X_6631_ la_data_in[20] _6631_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_20_614 VGND VPWR sky130_fd_sc_hd__decap_12
X_3843_ _3843_/A _4667_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_149_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_928 VGND VPWR sky130_fd_sc_hd__decap_12
X_3774_ _3773_/X _3767_/B _3774_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_6562_ _6495_/A la_data_in[13] _6497_/X _6562_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_121_1011 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_146_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_164_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_5513_ _5506_/X _5508_/X _5505_/X _5509_/X _5513_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_160_1093 VGND VPWR sky130_fd_sc_hd__decap_12
X_6493_ la_data_in[14] _6493_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_145_365 VGND VPWR sky130_fd_sc_hd__fill_1
X_5444_ _5444_/A _5444_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_121_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_1156 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_201_1090 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_145_398 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_160_335 VGND VPWR sky130_fd_sc_hd__fill_1
X_5375_ _5353_/X _5354_/X _5352_/X _5355_/X _5375_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_99_452 VGND VPWR sky130_fd_sc_hd__decap_12
X_7114_ _6905_/A _7114_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_4326_ _4272_/X _4273_/X _4272_/X _4273_/X _4326_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_102_947 VGND VPWR sky130_fd_sc_hd__decap_12
X_4257_ _4233_/X _4243_/X _4233_/X _4243_/X _4257_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_7045_ _7043_/Y _7044_/Y _7045_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_101_457 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_703 VGND VPWR sky130_fd_sc_hd__decap_12
X_4188_ _3693_/X _4235_/B _4190_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_132_1162 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_360 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_419 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_82_374 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_227 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_208_1222 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_179_27 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_452 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6829_ la_data_in[59] _6830_/B VGND VPWR sky130_fd_sc_hd__inv_8
XPHY_2259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_446 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_102 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_608 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_1130 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_195_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_630 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_136_321 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_1147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_195_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_855 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_1128 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_192_983 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_505 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_164_696 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_136_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_163_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_357 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_560 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_700 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_625 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_378 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_389 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_617 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_799 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_382 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_864 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_886 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_739 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_216 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_780 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_964 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_202_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_1011 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_187_733 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_148_1191 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_183_1082 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_175_928 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_293 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_186_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_822 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_146_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_833 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_1258 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_877 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_640 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_313 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_170_666 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_912 VGND VPWR sky130_fd_sc_hd__decap_3
X_5160_ _5155_/X _5159_/X _5158_/X _5160_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_111_700 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_571 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_1045 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_422 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_636 VGND VPWR sky130_fd_sc_hd__decap_12
X_4111_ _4089_/X _4090_/X _4089_/X _4090_/X _4111_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_155_1184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_733 VGND VPWR sky130_fd_sc_hd__decap_8
X_5091_ _5077_/X _5083_/X _5089_/X _5090_/X _5091_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_96_455 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_97_989 VGND VPWR sky130_fd_sc_hd__decap_12
X_4042_ _5294_/A _3933_/X _4044_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_204_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_522 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_209_152 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_864 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_209_196 VGND VPWR sky130_fd_sc_hd__decap_6
X_7801_ _3849_/Y _3842_/A _7801_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_363 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_823 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_92_694 VGND VPWR sky130_fd_sc_hd__decap_8
X_5993_ _5724_/X _5766_/X _5993_/C _5993_/D _5993_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_91_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_227 VGND VPWR sky130_fd_sc_hd__decap_12
X_7732_ _7732_/D _4475_/A _7801_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4944_ _4941_/X _4942_/X _4941_/X _4942_/X _4944_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_205_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_1005 VGND VPWR sky130_fd_sc_hd__decap_12
X_7663_ _6890_/X _6822_/A _7624_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_178_755 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_794 VGND VPWR sky130_fd_sc_hd__decap_12
X_4875_ _4675_/X _4689_/X _4622_/X _4690_/X _4875_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_177_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_1106 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_271 VGND VPWR sky130_fd_sc_hd__decap_4
X_6614_ _6612_/Y _6613_/Y _6614_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_178_788 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_800 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_20_444 VGND VPWR sky130_fd_sc_hd__decap_12
X_3826_ _3826_/A _4453_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_7594_ _7594_/HI la_data_out[121] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_192_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_989 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_758 VGND VPWR sky130_fd_sc_hd__decap_12
X_6545_ _6545_/A _6544_/X _6545_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_3757_ _3757_/A _3767_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_180_408 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_1196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_146_663 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_174_983 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_888 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_825 VGND VPWR sky130_fd_sc_hd__decap_3
X_6476_ _6466_/X _6476_/B _6475_/Y _7719_/D VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_161_611 VGND VPWR sky130_fd_sc_hd__decap_12
X_3688_ _6190_/A _3733_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_145_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_847 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_1191 VGND VPWR sky130_fd_sc_hd__decap_12
X_5427_ _5162_/A _4562_/B _5427_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_47_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_160_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_805 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_379 VGND VPWR sky130_fd_sc_hd__fill_1
X_5358_ _5338_/X _5346_/X _5356_/X _5357_/X _5358_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_102_711 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_838 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_593 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_293 VGND VPWR sky130_fd_sc_hd__decap_12
X_4309_ _4309_/A _4303_/X _4309_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_59_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_1129 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_181_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_232 VGND VPWR sky130_fd_sc_hd__decap_12
X_5289_ _5071_/X _5118_/X _5061_/X _5119_/X _5289_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_59_168 VGND VPWR sky130_fd_sc_hd__decap_12
X_7028_ _6970_/X _7027_/X _7024_/X _7028_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_74_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_190 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_210_1178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_739 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_1006 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_167_1077 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_867 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_167_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_1203 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_761 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_169_733 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_142_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_184_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_1217 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_293 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_2089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_168_276 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_196_596 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_415 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_74 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_104_1050 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_183_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_139_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_343 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_696 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_151_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_1184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_709 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_155_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_140_817 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_155_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_839 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_891 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_444 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_959 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_609 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_1054 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_812 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_206_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_344 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_569 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_159_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_794 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_3291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_43 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_175_703 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_202_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_574 VGND VPWR sky130_fd_sc_hd__decap_12
X_4660_ _4653_/X _4659_/X _4658_/X _4660_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_174_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_764 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_2590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_797 VGND VPWR sky130_fd_sc_hd__decap_6
X_4591_ _4547_/A _4591_/B _4592_/B VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_196_80 VGND VPWR sky130_fd_sc_hd__decap_12
X_6330_ _3933_/X _6334_/B _6332_/B VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_190_728 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_143_600 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_128_674 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_143_611 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_825 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_1077 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_696 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_1099 VGND VPWR sky130_fd_sc_hd__decap_12
X_6261_ _5724_/X _6260_/Y _6261_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_116_869 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_709 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_171_975 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_115_357 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_157_1257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_508 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_154 VGND VPWR sky130_fd_sc_hd__decap_12
X_5212_ _5207_/X _5208_/X _5207_/X _5208_/X _5212_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_130_316 VGND VPWR sky130_fd_sc_hd__decap_12
X_6192_ _6192_/A _6191_/X _7771_/D VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_170_496 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_349 VGND VPWR sky130_fd_sc_hd__decap_12
X_5143_ _4653_/A _4847_/B _5143_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_9_1056 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_477 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_263 VGND VPWR sky130_fd_sc_hd__decap_12
X_5074_ _4718_/A _4625_/B _5074_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4025_ _4005_/X _4023_/X _4021_/X _4024_/X _4025_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_37_330 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_491 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_839 VGND VPWR sky130_fd_sc_hd__decap_12
X_5976_ _5955_/X _5961_/X _5963_/X _5977_/B VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_164_1239 VGND VPWR sky130_fd_sc_hd__decap_12
X_7715_ _6488_/X _6421_/A _7785_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_4927_ _4926_/A _4926_/B _4926_/X _4927_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_21_731 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_166_703 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_178_563 VGND VPWR sky130_fd_sc_hd__decap_12
X_7646_ _7646_/D _6932_/A _7754_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_100_68 VGND VPWR sky130_fd_sc_hd__decap_12
X_4858_ _4857_/A _4856_/X _4857_/X _4858_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_166_736 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_205_1269 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_28 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_193_544 VGND VPWR sky130_fd_sc_hd__decap_4
X_3809_ _3791_/A _3807_/X _3808_/Y _3809_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_7577_ _7577_/HI la_data_out[104] VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_197_1026 VGND VPWR sky130_fd_sc_hd__decap_8
X_4789_ _4785_/X _4788_/X _4785_/X _4788_/X _4789_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_165_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_652 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_419 VGND VPWR sky130_fd_sc_hd__decap_8
X_6528_ _7700_/Q _6530_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_146_471 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_101_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_180_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_1139 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_6459_ _6439_/X _6458_/X _6455_/X _6459_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_161_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_192_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_602 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_891 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_1062 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_850 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_764 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_872 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_1065 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_134_1076 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_894 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_425 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_959 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_1240 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_1202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_853 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_169_1128 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_875 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_812 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_85 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_189_806 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_141 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_188_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_203_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_1060 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_697 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_388 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_1191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_51 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_157_714 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_230 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_156_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_764 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_211_180 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_141_1036 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_200_898 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_156_279 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_61 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_994 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_941 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_153_964 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_655 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_828 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_1151 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_112_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_904 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_775 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_756 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_187_1217 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_943 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_428 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_207_464 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_322 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_642 VGND VPWR sky130_fd_sc_hd__decap_12
X_5830_ _5826_/X _5829_/X _5826_/X _5829_/X _5830_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_90_973 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_675 VGND VPWR sky130_fd_sc_hd__decap_12
X_5761_ _5726_/X _5759_/X _5726_/X _5759_/X _5761_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_210_629 VGND VPWR sky130_fd_sc_hd__decap_12
X_7500_ _7500_/HI la_data_out[27] VGND VPWR sky130_fd_sc_hd__conb_1
X_4712_ _4707_/X _4708_/X _4707_/X _4708_/X _4712_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_188_883 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_1166 VGND VPWR sky130_fd_sc_hd__decap_12
X_5692_ _5690_/X _5691_/X _5692_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_72_1199 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_30_572 VGND VPWR sky130_fd_sc_hd__decap_8
X_7431_ io_oeb[26] _7431_/LO VGND VPWR sky130_fd_sc_hd__conb_1
X_4643_ _4642_/A _4642_/B _4642_/X _4643_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_175_566 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_717 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_419 VGND VPWR sky130_fd_sc_hd__decap_8
X_7362_ _5059_/Y _7355_/X _7361_/X wbs_dat_o[17] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_116_611 VGND VPWR sky130_fd_sc_hd__decap_12
X_4574_ _4497_/X _4501_/X _4500_/X _4574_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_162_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_471 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_1166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_110 VGND VPWR sky130_fd_sc_hd__decap_12
X_6313_ _5972_/A _5972_/B _5973_/X _6313_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_157_1021 VGND VPWR sky130_fd_sc_hd__decap_12
X_7293_ _7370_/A _7293_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_131_603 VGND VPWR sky130_fd_sc_hd__decap_6
X_6244_ _5277_/Y _6216_/X _6194_/X _6244_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_171_794 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_157_1087 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_29 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_658 VGND VPWR sky130_fd_sc_hd__decap_12
X_6175_ _6151_/X _6176_/B VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_97_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_712 VGND VPWR sky130_fd_sc_hd__decap_12
X_5126_ _5125_/A _5125_/B _5125_/X _5126_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_97_594 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_745 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_959 VGND VPWR sky130_fd_sc_hd__decap_12
X_5057_ _5055_/X _5056_/X _5054_/X _5057_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XPHY_4706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4008_ _4568_/A _3949_/B _4008_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_84_288 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_845 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_1123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_197_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_483 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_1099 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_27 VGND VPWR sky130_fd_sc_hd__decap_12
X_5959_ _5932_/X _5933_/X _5934_/X _5959_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_164_1069 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_200_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_187_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_1206 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_550 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_583 VGND VPWR sky130_fd_sc_hd__decap_12
X_7629_ _7629_/D _7043_/A _7729_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_193_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_205_1099 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_886 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_181_525 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_780 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_611 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_1162 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_964 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_162_761 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_1135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_1105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_883 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_723 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_948 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_487 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_691 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_95 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_789 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_428 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_1111 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_1182 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_620 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_642 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_189_625 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_204_434 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_1117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_889 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_147_1245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_1008 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_837 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_483 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_350 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_361 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_372 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_383 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_157_522 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_185_842 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_394 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_196_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_565 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_184_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_144_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_4 _4498_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_290 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_1221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_153_761 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_1257 VGND VPWR sky130_fd_sc_hd__decap_12
X_4290_ _4289_/Y _4291_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_153_794 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_496 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_636 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_369 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_403 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_1004 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_1082 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_745 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_767 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_929 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_575 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_208_740 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_417 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_981 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_288 VGND VPWR sky130_fd_sc_hd__decap_12
X_6931_ _6929_/Y _6931_/B _6931_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_187_1069 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_208_784 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_951 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_208_795 VGND VPWR sky130_fd_sc_hd__decap_12
X_6862_ _6922_/A _6861_/X _6862_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_81_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_303 VGND VPWR sky130_fd_sc_hd__decap_12
X_5813_ _5803_/X _5804_/X _5803_/X _5804_/X _5813_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_179_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_483 VGND VPWR sky130_fd_sc_hd__decap_12
X_6793_ _6795_/A _6764_/X _6792_/Y _6793_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_204_990 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_194_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_1061 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_358 VGND VPWR sky130_fd_sc_hd__decap_4
X_5744_ _5729_/X _5735_/X _5742_/X _5743_/X _5745_/B VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_148_511 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_148_544 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_864 VGND VPWR sky130_fd_sc_hd__decap_12
X_5675_ _5665_/X _5672_/X _5673_/X _5674_/X _5675_/X VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_202_1239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_886 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_191_812 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_1086 VGND VPWR sky130_fd_sc_hd__decap_12
X_7414_ io_oeb[9] _7414_/LO VGND VPWR sky130_fd_sc_hd__conb_1
XFILLER_190_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_1154 VGND VPWR sky130_fd_sc_hd__decap_12
X_4626_ _3811_/A _5095_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_191_834 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_547 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_191_867 VGND VPWR sky130_fd_sc_hd__decap_12
X_7345_ _7345_/A _7351_/B _7345_/X VGND VPWR sky130_fd_sc_hd__or2_4
X_4557_ _4552_/X _4556_/X _4552_/X _4556_/X _4557_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_144_772 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_934 VGND VPWR sky130_fd_sc_hd__decap_12
X_7276_ _7276_/A _7300_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_104_636 VGND VPWR sky130_fd_sc_hd__decap_4
X_4488_ _7731_/Q _4488_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_103_135 VGND VPWR sky130_fd_sc_hd__decap_12
X_6227_ _6228_/A _6228_/B _6227_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_135_1160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_56 VGND VPWR sky130_fd_sc_hd__decap_12
X_6158_ _6158_/A _6158_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_66_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_391 VGND VPWR sky130_fd_sc_hd__decap_12
X_5109_ _4548_/A _4505_/B _5111_/A VGND VPWR sky130_fd_sc_hd__or2_4
X_6089_ _6219_/A _6089_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_100_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_1139 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_428 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_17_119 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_4503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_122_44 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_759 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_491 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_4536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_642 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_4547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_4569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_198_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_198_422 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_623 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_837 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_3868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_3879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_201_415 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_1101 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_318 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_1003 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_1183 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_142_1142 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_178_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_210_971 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_1156 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_166_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_193_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_513 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_182_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_147_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_452 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_912 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_422 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_150_753 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_730 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_150_764 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_818 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_1_752 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_606 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_150_786 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_163_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_892 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_520 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_1266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_778 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_501 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_726 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_82 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_93 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_940 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_483 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_1015 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_943 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_60_965 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_176_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_807 VGND VPWR sky130_fd_sc_hd__decap_12
X_3790_ wbs_dat_i[14] _3790_/B _3790_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_31_166 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_180 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_191 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_160_1264 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_158_886 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_185_672 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_172_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_739 VGND VPWR sky130_fd_sc_hd__decap_12
X_5460_ _5455_/X _5458_/A _5459_/X _6198_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_68_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_173_867 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_145_558 VGND VPWR sky130_fd_sc_hd__decap_3
X_4411_ _4409_/X _4410_/X _4408_/X _4411_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_5391_ _5336_/X _5380_/X _5389_/X _5390_/X _5391_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_7130_ _7128_/A _7130_/B _7129_/Y _7130_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_4342_ _4919_/A _4461_/B _4342_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_158_1171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_945 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_153_591 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_141_753 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_807 VGND VPWR sky130_fd_sc_hd__decap_12
X_7061_ _7623_/Q _7061_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_193_1095 VGND VPWR sky130_fd_sc_hd__decap_3
X_4273_ _4259_/X _4266_/X _4259_/X _4266_/X _4273_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_154_1057 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_141_786 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_140_263 VGND VPWR sky130_fd_sc_hd__decap_12
X_6012_ _4991_/X _6012_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_100_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_499 VGND VPWR sky130_fd_sc_hd__decap_12
.ends

