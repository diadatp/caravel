magic
tech sky130A
magscale 1 2
timestamp 1607074398
<< checkpaint >>
rect -9696 -8626 593620 712562
<< locali >>
rect 154313 676243 154347 685797
rect 218989 666587 219023 676141
rect 494069 666587 494103 676141
rect 542737 666587 542771 684437
rect 559297 666587 559331 684437
rect 219265 647275 219299 656829
rect 219357 616879 219391 626501
rect 219081 608719 219115 611405
rect 219265 601579 219299 608549
rect 542553 601715 542587 608549
rect 559113 601715 559147 608549
rect 219173 589339 219207 598893
rect 542737 589339 542771 598893
rect 559297 589339 559331 598893
rect 154313 579751 154347 589237
rect 218897 569959 218931 579581
rect 494161 563091 494195 569857
rect 218897 550647 218931 553401
rect 542461 550647 542495 560201
rect 559021 550647 559055 560201
rect 154405 521679 154439 531233
rect 154405 502367 154439 511921
rect 219081 505087 219115 510561
rect 542553 485775 542587 492609
rect 559113 485775 559147 492609
rect 154405 476051 154439 482953
rect 542553 463743 542587 466497
rect 559113 463743 559147 466497
rect 96629 463267 96663 463369
rect 89729 463131 89763 463233
rect 106197 463199 106231 463369
rect 125609 463199 125643 463301
rect 157349 463131 157383 463369
rect 160937 463267 160971 463369
rect 118651 463097 118709 463131
rect 173909 462995 173943 463233
rect 183569 463199 183603 463369
rect 193137 463199 193171 463369
rect 195897 463199 195931 463233
rect 195839 463165 195931 463199
rect 200129 463199 200163 463369
rect 205649 463199 205683 463369
rect 259469 463199 259503 463505
rect 222243 463165 222301 463199
rect 234571 463165 234629 463199
rect 244231 463165 244289 463199
rect 253891 463165 253949 463199
rect 269037 463199 269071 463505
rect 269129 463267 269163 463505
rect 278697 463267 278731 463505
rect 282929 463403 282963 463573
rect 286977 463471 287011 463641
rect 287069 463471 287103 463505
rect 287069 463437 287253 463471
rect 287713 463403 287747 463505
rect 283021 463267 283055 463369
rect 287805 463267 287839 463573
rect 291209 463199 291243 463437
rect 291301 463267 291335 463437
rect 293601 463335 293635 463573
rect 296637 463267 296671 463505
rect 183477 462995 183511 463165
rect 280019 463029 280261 463063
rect 6929 459119 6963 459425
rect 16497 459255 16531 459425
rect 16589 459119 16623 459221
rect 26249 459119 26283 459425
rect 35817 459255 35851 459425
rect 35909 459119 35943 459221
rect 45569 459119 45603 459425
rect 55137 459255 55171 459425
rect 55229 459119 55263 459221
rect 64889 459119 64923 459425
rect 74457 459255 74491 459425
rect 74549 459119 74583 459221
rect 84853 459119 84887 459425
rect 94513 459119 94547 459425
rect 104173 459119 104207 459425
rect 113833 459119 113867 459425
rect 123493 459119 123527 459425
rect 133153 459119 133187 459425
rect 142813 459119 142847 459425
rect 152473 459119 152507 459425
rect 162133 459119 162167 459425
rect 171793 459119 171827 459425
rect 181453 459119 181487 459425
rect 191113 459119 191147 459425
rect 200773 459119 200807 459425
rect 210433 459119 210467 459425
rect 220093 459119 220127 459425
rect 225337 459119 225371 459425
rect 234629 459119 234663 459221
rect 238033 458235 238067 459425
rect 240057 458303 240091 459425
rect 243369 458507 243403 459425
rect 246497 458575 246531 459425
rect 247417 459255 247451 459493
rect 249625 458847 249659 459425
rect 254961 459119 254995 459425
rect 258733 459255 258767 459493
rect 268393 459255 268427 459493
rect 278053 459255 278087 459493
rect 287713 459255 287747 459493
rect 296637 459255 296671 459493
rect 306389 459255 306423 459493
rect 315957 459255 315991 459493
rect 331229 458983 331263 459289
rect 332149 459051 332183 459289
rect 334173 458915 334207 459289
rect 335369 458779 335403 459289
rect 337301 458711 337335 459289
rect 338405 458643 338439 459289
rect 340705 458439 340739 459289
rect 341533 458371 341567 459289
rect 317889 338147 317923 340153
rect 326261 337501 326445 337535
rect 326261 337467 326295 337501
rect 331137 336719 331171 337433
rect 100677 318835 100711 328389
rect 107485 327131 107519 336685
rect 331229 336719 331263 337433
rect 232145 328491 232179 335733
rect 244473 328491 244507 334441
rect 231133 318835 231167 328389
rect 254685 318835 254719 328389
rect 257077 317475 257111 327029
rect 262781 325703 262815 333693
rect 279525 327131 279559 336685
rect 280629 318835 280663 328389
rect 281917 318835 281951 328389
rect 295625 322235 295659 327029
rect 319453 325703 319487 328389
rect 320281 325703 320315 335189
rect 100677 299523 100711 309077
rect 107485 307819 107519 317373
rect 244381 311491 244415 317373
rect 238033 299523 238067 309077
rect 100677 280211 100711 289765
rect 107485 288439 107519 298061
rect 231225 289867 231259 299421
rect 232421 288439 232455 298061
rect 240701 289867 240735 299421
rect 238033 280211 238067 289765
rect 231225 270555 231259 280109
rect 240701 270555 240735 280109
rect 245025 278783 245059 298061
rect 257077 294491 257111 302889
rect 258825 298163 258859 315945
rect 260389 307819 260423 317373
rect 261585 299523 261619 317373
rect 265817 307887 265851 317373
rect 282653 309179 282687 318665
rect 335829 316047 335863 325601
rect 341625 317475 341659 327029
rect 344293 318835 344327 328389
rect 260297 289867 260331 299421
rect 264529 298163 264563 307717
rect 265817 298163 265851 307717
rect 293417 306391 293451 309145
rect 316877 298163 316911 307717
rect 319453 306391 319487 315945
rect 320281 306391 320315 315945
rect 339969 307819 340003 317373
rect 246037 270555 246071 280109
rect 246405 278783 246439 288337
rect 257169 278783 257203 280109
rect 258733 277423 258767 286977
rect 265817 278851 265851 288337
rect 319637 287079 319671 298061
rect 321109 288507 321143 298061
rect 333161 288439 333195 289969
rect 339969 282863 340003 298061
rect 100677 260899 100711 270453
rect 238033 260899 238067 270453
rect 260297 265319 260331 273241
rect 264529 269127 264563 278681
rect 265817 269127 265851 278681
rect 231225 251243 231259 260797
rect 322305 259471 322339 263585
rect 232145 253895 232179 258009
rect 232421 253215 232455 258009
rect 100677 241519 100711 251141
rect 244381 241587 244415 258009
rect 256985 249815 257019 251209
rect 232697 235331 232731 240057
rect 246313 238799 246347 248353
rect 258825 240227 258859 249713
rect 299029 247095 299063 256649
rect 232053 230503 232087 234617
rect 261585 234583 261619 238697
rect 300317 237439 300351 246993
rect 301789 237439 301823 246993
rect 319637 240159 319671 258009
rect 326261 249815 326295 254065
rect 334541 251107 334575 256649
rect 335737 250971 335771 258009
rect 341625 251243 341659 260797
rect 232053 222207 232087 224961
rect 260389 224247 260423 229041
rect 299029 227783 299063 237337
rect 246405 209831 246439 217413
rect 260389 214523 260423 219385
rect 261585 215271 261619 219385
rect 299029 218059 299063 227613
rect 300317 218059 300351 227681
rect 301789 226355 301823 235909
rect 330401 230095 330435 235909
rect 244473 201535 244507 202861
rect 300317 198747 300351 208301
rect 301789 207043 301823 216597
rect 319637 209831 319671 219385
rect 321109 209831 321143 219385
rect 322121 209831 322155 219317
rect 333069 218059 333103 227681
rect 340061 220779 340095 229041
rect 326261 200175 326295 215373
rect 329021 205683 329055 215237
rect 334633 207043 334667 216597
rect 232329 172567 232363 182121
rect 244381 173927 244415 189465
rect 244933 183583 244967 195245
rect 260205 183515 260239 191777
rect 261493 182155 261527 190417
rect 260297 173859 260331 182121
rect 263057 180863 263091 190417
rect 299029 189091 299063 198645
rect 264529 171139 264563 180761
rect 265817 171139 265851 180761
rect 293141 171139 293175 180761
rect 300317 179435 300351 188989
rect 301789 187731 301823 197149
rect 319637 190519 319671 200073
rect 321109 190519 321143 200073
rect 322213 190519 322247 200073
rect 329021 187731 329055 197285
rect 330585 187731 330619 205581
rect 335829 203575 335863 209729
rect 340061 204935 340095 211089
rect 334633 187731 334667 197285
rect 333161 182087 333195 183889
rect 335829 180863 335863 190417
rect 107485 153255 107519 162809
rect 232605 153187 232639 161381
rect 232053 143599 232087 153153
rect 253029 151827 253063 161381
rect 257077 151827 257111 161381
rect 107485 133943 107519 143497
rect 231225 135371 231259 137989
rect 232053 132515 232087 142069
rect 100677 106335 100711 115889
rect 107485 114563 107519 124117
rect 232421 118711 232455 136425
rect 240701 133943 240735 143497
rect 244933 131223 244967 140709
rect 246037 133331 246071 143497
rect 246405 142171 246439 143565
rect 253029 142239 253063 151657
rect 260297 149107 260331 158661
rect 293325 151827 293359 161381
rect 299029 160123 299063 169677
rect 300317 160123 300351 169677
rect 301789 168419 301823 177973
rect 319637 171139 319671 180761
rect 321109 171139 321143 180761
rect 334541 179503 334575 180829
rect 334541 171071 334575 179333
rect 319637 151827 319671 161381
rect 321109 151827 321143 161381
rect 326353 161347 326387 169677
rect 331781 168419 331815 169813
rect 246405 124219 246439 141865
rect 253213 131155 253247 140709
rect 258825 138635 258859 143497
rect 264529 142171 264563 151725
rect 260205 129795 260239 139349
rect 293325 132515 293359 142069
rect 296085 140811 296119 150365
rect 301513 147679 301547 150229
rect 231225 116059 231259 118677
rect 231225 106335 231259 115889
rect 244381 113203 244415 122757
rect 245025 113135 245059 121397
rect 100677 87023 100711 96577
rect 107485 95251 107519 104805
rect 231225 96747 231259 99365
rect 232145 92531 232179 102085
rect 232329 93891 232363 106981
rect 244381 103615 244415 113033
rect 253121 108375 253155 122757
rect 254685 104907 254719 122757
rect 257169 113203 257203 122757
rect 261493 122723 261527 131053
rect 299029 129863 299063 140709
rect 300317 130747 300351 140709
rect 301881 140675 301915 141049
rect 314393 138499 314427 143497
rect 258917 106335 258951 115889
rect 260389 106335 260423 115889
rect 261493 111843 261527 121261
rect 263057 104907 263091 117997
rect 264621 113203 264655 122757
rect 265817 113203 265851 122757
rect 299029 120207 299063 129693
rect 301789 121499 301823 134521
rect 319637 132515 319671 142069
rect 330493 140811 330527 150365
rect 331781 142171 331815 151725
rect 334541 142171 334575 151725
rect 329021 131155 329055 140709
rect 331781 131155 331815 140709
rect 335921 131155 335955 140709
rect 294797 103547 294831 113101
rect 246313 95183 246347 99433
rect 253213 95183 253247 103445
rect 100677 67643 100711 77197
rect 107485 75939 107519 85493
rect 232329 75939 232363 89709
rect 253029 84235 253063 85629
rect 257077 85595 257111 95149
rect 258917 93891 258951 103445
rect 261585 85527 261619 99773
rect 263057 93891 263091 103445
rect 264437 93891 264471 103445
rect 265725 95183 265759 103445
rect 293325 93891 293359 103445
rect 297465 100759 297499 106913
rect 298937 102187 298971 120037
rect 300225 102187 300259 120037
rect 301697 102187 301731 120037
rect 317153 117555 317187 124117
rect 317337 115583 317371 124117
rect 316969 104907 317003 114461
rect 317153 107627 317187 114461
rect 317245 106131 317279 114393
rect 317337 109735 317371 114461
rect 319637 113203 319671 122621
rect 334449 121499 334483 131053
rect 340061 124219 340095 133841
rect 319637 93891 319671 103445
rect 321109 93891 321143 106029
rect 326169 103547 326203 113101
rect 331781 111843 331815 121397
rect 322305 93891 322339 103445
rect 334541 102255 334575 111741
rect 335829 103615 335863 113101
rect 339969 108987 340003 115481
rect 328929 92531 328963 102085
rect 334541 92531 334575 102085
rect 335921 93891 335955 103445
rect 296637 86887 296671 89029
rect 340061 85595 340095 95149
rect 244473 77231 244507 84133
rect 246037 74579 246071 77333
rect 100677 48331 100711 57885
rect 107485 56627 107519 66181
rect 100677 29019 100711 38573
rect 107485 37315 107519 46869
rect 231317 45611 231351 55165
rect 232145 46971 232179 73049
rect 253213 63563 253247 73117
rect 254777 69683 254811 75837
rect 261677 74647 261711 84133
rect 263057 67643 263091 82977
rect 264529 74579 264563 84133
rect 293325 74579 293359 84133
rect 294797 74579 294831 84133
rect 314209 67643 314243 77197
rect 318165 67643 318199 77197
rect 319637 74579 319671 84133
rect 320833 82943 320867 84269
rect 320833 73219 320867 82773
rect 329021 71791 329055 82773
rect 240609 47039 240643 56525
rect 244473 46971 244507 56525
rect 246497 48331 246531 57885
rect 254777 53839 254811 63461
rect 261585 46971 261619 55981
rect 264529 46971 264563 64821
rect 265817 55335 265851 64821
rect 232329 27659 232363 40681
rect 232789 27659 232823 40681
rect 240701 37383 240735 46869
rect 265817 45611 265851 55165
rect 293325 46971 293359 64821
rect 294797 46971 294831 64821
rect 296085 46971 296119 59993
rect 314209 56627 314243 66181
rect 299029 45611 299063 55165
rect 300317 45611 300351 55165
rect 301789 45611 301823 55165
rect 319637 46971 319671 64821
rect 244381 38607 244415 41429
rect 252937 40715 252971 45509
rect 107485 9707 107519 27557
rect 244473 18003 244507 27557
rect 252937 26299 252971 35853
rect 257169 27659 257203 45509
rect 261585 35955 261619 42109
rect 264437 35955 264471 45509
rect 265725 35955 265759 37349
rect 314209 37315 314243 46869
rect 321017 45611 321051 63461
rect 322305 55335 322339 64821
rect 331781 53839 331815 63461
rect 334541 46971 334575 61421
rect 345397 57987 345431 67541
rect 319637 35955 319671 45509
rect 322305 40715 322339 45509
rect 299029 26299 299063 35853
rect 300317 26299 300351 35853
rect 301789 26299 301823 35853
rect 321017 31739 321051 40681
rect 326353 27659 326387 44081
rect 231133 16507 231167 16541
rect 231317 16541 231409 16575
rect 231317 16507 231351 16541
rect 231133 16473 231351 16507
rect 268761 13107 268795 16677
rect 268853 12563 268887 16609
rect 268945 13175 268979 16677
rect 269037 13107 269071 16609
rect 278237 12767 278271 17085
rect 278329 12835 278363 17085
rect 278421 9639 278455 17153
rect 55263 3825 55447 3859
rect 55263 3689 55355 3723
rect 34621 3383 34655 3621
rect 55229 3315 55263 3553
rect 55321 3247 55355 3689
rect 55413 3179 55447 3825
rect 58725 3383 58759 4097
rect 64521 3825 64797 3859
rect 64521 3179 64555 3825
rect 64613 3689 64797 3723
rect 64613 3247 64647 3689
rect 64797 3315 64831 3553
rect 64739 3281 64831 3315
rect 64889 3179 64923 3621
rect 74457 3179 74491 3621
rect 84209 3043 84243 3621
rect 90925 595 90959 9605
rect 99297 2975 99331 3621
rect 100493 595 100527 9605
rect 101505 2839 101539 3621
rect 108773 595 108807 9605
rect 278513 9571 278547 17085
rect 278605 12087 278639 17153
rect 278697 13107 278731 17085
rect 297557 13991 297591 23341
rect 300685 14059 300719 23409
rect 301789 14399 301823 18241
rect 301881 14331 301915 18173
rect 301973 15215 302007 17221
rect 302065 15147 302099 17289
rect 302157 15215 302191 17221
rect 304641 15215 304675 18037
rect 314209 18003 314243 27557
rect 304917 15215 304951 17969
rect 329113 15215 329147 17969
rect 307217 11407 307251 15181
rect 322673 9129 323133 9163
rect 322673 9095 322707 9129
rect 322765 9061 323041 9095
rect 322765 9027 322799 9061
rect 324053 8993 324513 9027
rect 324053 8959 324087 8993
rect 345397 8347 345431 11033
rect 135303 4709 135453 4743
rect 154623 4709 154773 4743
rect 125609 4471 125643 4573
rect 135177 4471 135211 4641
rect 135361 4539 135395 4641
rect 144929 4403 144963 4505
rect 154497 4403 154531 4641
rect 154589 4403 154623 4573
rect 238769 4539 238803 4573
rect 239413 4573 239689 4607
rect 239413 4539 239447 4573
rect 238769 4505 239045 4539
rect 164157 4403 164191 4505
rect 246681 4471 246715 4573
rect 250269 4471 250303 5525
rect 252937 5423 252971 8245
rect 267289 5355 267323 5525
rect 268393 5355 268427 5525
rect 268301 4947 268335 5321
rect 263425 4403 263459 4505
rect 264989 4403 265023 4777
rect 267381 4335 267415 4845
rect 270693 4743 270727 5049
rect 128277 3655 128311 4165
rect 117053 3621 117329 3655
rect 117053 2839 117087 3621
rect 119353 2975 119387 3621
rect 128369 3655 128403 4165
rect 147597 3655 147631 4165
rect 157257 3655 157291 4165
rect 168665 3893 168883 3927
rect 124229 3043 124263 3621
rect 168665 3587 168699 3893
rect 168849 3859 168883 3893
rect 171701 3893 171919 3927
rect 171701 3859 171735 3893
rect 168757 3587 168791 3825
rect 171793 3655 171827 3825
rect 171885 3383 171919 3893
rect 171793 3315 171827 3349
rect 171977 3315 172011 3689
rect 176485 3383 176519 4165
rect 176577 3655 176611 4301
rect 180533 3383 180567 3689
rect 180625 3587 180659 3825
rect 180717 3587 180751 4165
rect 180809 3655 180843 4165
rect 190377 3655 190411 4165
rect 200129 3655 200163 4165
rect 205741 3723 205775 4165
rect 180533 3349 180717 3383
rect 171793 3281 172011 3315
rect 208041 3315 208075 3553
rect 208133 3383 208167 3553
rect 215033 3383 215067 4165
rect 215125 3655 215159 4301
rect 215217 3859 215251 4233
rect 215309 3859 215343 4233
rect 215401 3723 215435 4165
rect 215493 3383 215527 4301
rect 239229 4301 239505 4335
rect 264839 4301 265081 4335
rect 239229 4199 239263 4301
rect 268393 4267 268427 4709
rect 220185 3723 220219 4165
rect 270785 4199 270819 4709
rect 220093 3383 220127 3553
rect 208225 3315 208259 3349
rect 208041 3281 208259 3315
rect 220001 3315 220035 3349
rect 220277 3315 220311 3689
rect 224877 3587 224911 4165
rect 263643 3825 263735 3859
rect 263701 3587 263735 3825
rect 220001 3281 220311 3315
rect 266001 3315 266035 3553
rect 266093 3383 266127 3553
rect 270509 3383 270543 3621
rect 277961 3621 278179 3655
rect 277961 3383 277995 3621
rect 278145 3587 278179 3621
rect 266185 3315 266219 3349
rect 266001 3281 266219 3315
rect 278053 3383 278087 3553
rect 124137 3009 124263 3043
rect 124137 2975 124171 3009
rect 124229 2771 124263 2941
rect 267749 2771 267783 3349
rect 277317 2771 277351 3349
rect 280077 595 280111 6341
rect 282745 3859 282779 4233
rect 282837 3587 282871 3825
rect 282779 3553 282871 3587
rect 285321 3621 285539 3655
rect 285321 3587 285355 3621
rect 285413 3383 285447 3553
rect 285505 3383 285539 3621
rect 292405 3383 292439 4233
rect 292497 3859 292531 4301
rect 292589 3859 292623 4301
rect 292681 3383 292715 4233
rect 303813 3893 304123 3927
rect 303813 3723 303847 3893
rect 304089 3859 304123 3893
rect 306941 3893 307159 3927
rect 306941 3859 306975 3893
rect 303905 3587 303939 3689
rect 297373 3383 297407 3553
rect 303997 3587 304031 3825
rect 297281 3315 297315 3349
rect 297465 3315 297499 3553
rect 297281 3281 297499 3315
rect 306849 3315 306883 3689
rect 306941 3383 306975 3689
rect 307033 3655 307067 3825
rect 307125 3655 307159 3893
rect 316693 3893 316911 3927
rect 316693 3859 316727 3893
rect 313657 3383 313691 3621
rect 313749 3383 313783 3689
rect 316785 3587 316819 3825
rect 316877 3655 316911 3893
rect 316877 3621 317061 3655
rect 324973 3519 325007 3689
rect 326537 3655 326571 4165
rect 326295 3621 326571 3655
rect 326629 3383 326663 3621
rect 307033 3315 307067 3349
rect 306849 3281 307067 3315
<< viali >>
rect 154313 685797 154347 685831
rect 154313 676209 154347 676243
rect 542737 684437 542771 684471
rect 218989 676141 219023 676175
rect 218989 666553 219023 666587
rect 494069 676141 494103 676175
rect 494069 666553 494103 666587
rect 542737 666553 542771 666587
rect 559297 684437 559331 684471
rect 559297 666553 559331 666587
rect 219265 656829 219299 656863
rect 219265 647241 219299 647275
rect 219357 626501 219391 626535
rect 219357 616845 219391 616879
rect 219081 611405 219115 611439
rect 219081 608685 219115 608719
rect 219265 608549 219299 608583
rect 542553 608549 542587 608583
rect 542553 601681 542587 601715
rect 559113 608549 559147 608583
rect 559113 601681 559147 601715
rect 219265 601545 219299 601579
rect 219173 598893 219207 598927
rect 219173 589305 219207 589339
rect 542737 598893 542771 598927
rect 542737 589305 542771 589339
rect 559297 598893 559331 598927
rect 559297 589305 559331 589339
rect 154313 589237 154347 589271
rect 154313 579717 154347 579751
rect 218897 579581 218931 579615
rect 218897 569925 218931 569959
rect 494161 569857 494195 569891
rect 494161 563057 494195 563091
rect 542461 560201 542495 560235
rect 218897 553401 218931 553435
rect 218897 550613 218931 550647
rect 542461 550613 542495 550647
rect 559021 560201 559055 560235
rect 559021 550613 559055 550647
rect 154405 531233 154439 531267
rect 154405 521645 154439 521679
rect 154405 511921 154439 511955
rect 219081 510561 219115 510595
rect 219081 505053 219115 505087
rect 154405 502333 154439 502367
rect 542553 492609 542587 492643
rect 542553 485741 542587 485775
rect 559113 492609 559147 492643
rect 559113 485741 559147 485775
rect 154405 482953 154439 482987
rect 154405 476017 154439 476051
rect 542553 466497 542587 466531
rect 542553 463709 542587 463743
rect 559113 466497 559147 466531
rect 559113 463709 559147 463743
rect 286977 463641 287011 463675
rect 282929 463573 282963 463607
rect 259469 463505 259503 463539
rect 96629 463369 96663 463403
rect 89729 463233 89763 463267
rect 96629 463233 96663 463267
rect 106197 463369 106231 463403
rect 157349 463369 157383 463403
rect 106197 463165 106231 463199
rect 125609 463301 125643 463335
rect 125609 463165 125643 463199
rect 160937 463369 160971 463403
rect 183569 463369 183603 463403
rect 160937 463233 160971 463267
rect 173909 463233 173943 463267
rect 89729 463097 89763 463131
rect 118617 463097 118651 463131
rect 118709 463097 118743 463131
rect 157349 463097 157383 463131
rect 173909 462961 173943 462995
rect 183477 463165 183511 463199
rect 183569 463165 183603 463199
rect 193137 463369 193171 463403
rect 200129 463369 200163 463403
rect 195897 463233 195931 463267
rect 193137 463165 193171 463199
rect 195805 463165 195839 463199
rect 200129 463165 200163 463199
rect 205649 463369 205683 463403
rect 205649 463165 205683 463199
rect 222209 463165 222243 463199
rect 222301 463165 222335 463199
rect 234537 463165 234571 463199
rect 234629 463165 234663 463199
rect 244197 463165 244231 463199
rect 244289 463165 244323 463199
rect 253857 463165 253891 463199
rect 253949 463165 253983 463199
rect 259469 463165 259503 463199
rect 269037 463505 269071 463539
rect 269129 463505 269163 463539
rect 269129 463233 269163 463267
rect 278697 463505 278731 463539
rect 287805 463573 287839 463607
rect 286977 463437 287011 463471
rect 287069 463505 287103 463539
rect 287713 463505 287747 463539
rect 287253 463437 287287 463471
rect 282929 463369 282963 463403
rect 283021 463369 283055 463403
rect 287713 463369 287747 463403
rect 278697 463233 278731 463267
rect 283021 463233 283055 463267
rect 293601 463573 293635 463607
rect 287805 463233 287839 463267
rect 291209 463437 291243 463471
rect 269037 463165 269071 463199
rect 291301 463437 291335 463471
rect 293601 463301 293635 463335
rect 296637 463505 296671 463539
rect 291301 463233 291335 463267
rect 296637 463233 296671 463267
rect 291209 463165 291243 463199
rect 279985 463029 280019 463063
rect 280261 463029 280295 463063
rect 183477 462961 183511 462995
rect 247417 459493 247451 459527
rect 6929 459425 6963 459459
rect 16497 459425 16531 459459
rect 26249 459425 26283 459459
rect 16497 459221 16531 459255
rect 16589 459221 16623 459255
rect 6929 459085 6963 459119
rect 16589 459085 16623 459119
rect 35817 459425 35851 459459
rect 45569 459425 45603 459459
rect 35817 459221 35851 459255
rect 35909 459221 35943 459255
rect 26249 459085 26283 459119
rect 35909 459085 35943 459119
rect 55137 459425 55171 459459
rect 64889 459425 64923 459459
rect 55137 459221 55171 459255
rect 55229 459221 55263 459255
rect 45569 459085 45603 459119
rect 55229 459085 55263 459119
rect 74457 459425 74491 459459
rect 84853 459425 84887 459459
rect 74457 459221 74491 459255
rect 74549 459221 74583 459255
rect 64889 459085 64923 459119
rect 74549 459085 74583 459119
rect 84853 459085 84887 459119
rect 94513 459425 94547 459459
rect 94513 459085 94547 459119
rect 104173 459425 104207 459459
rect 104173 459085 104207 459119
rect 113833 459425 113867 459459
rect 113833 459085 113867 459119
rect 123493 459425 123527 459459
rect 123493 459085 123527 459119
rect 133153 459425 133187 459459
rect 133153 459085 133187 459119
rect 142813 459425 142847 459459
rect 142813 459085 142847 459119
rect 152473 459425 152507 459459
rect 152473 459085 152507 459119
rect 162133 459425 162167 459459
rect 162133 459085 162167 459119
rect 171793 459425 171827 459459
rect 171793 459085 171827 459119
rect 181453 459425 181487 459459
rect 181453 459085 181487 459119
rect 191113 459425 191147 459459
rect 191113 459085 191147 459119
rect 200773 459425 200807 459459
rect 200773 459085 200807 459119
rect 210433 459425 210467 459459
rect 210433 459085 210467 459119
rect 220093 459425 220127 459459
rect 220093 459085 220127 459119
rect 225337 459425 225371 459459
rect 238033 459425 238067 459459
rect 225337 459085 225371 459119
rect 234629 459221 234663 459255
rect 234629 459085 234663 459119
rect 240057 459425 240091 459459
rect 243369 459425 243403 459459
rect 246497 459425 246531 459459
rect 258733 459493 258767 459527
rect 247417 459221 247451 459255
rect 249625 459425 249659 459459
rect 254961 459425 254995 459459
rect 258733 459221 258767 459255
rect 268393 459493 268427 459527
rect 268393 459221 268427 459255
rect 278053 459493 278087 459527
rect 278053 459221 278087 459255
rect 287713 459493 287747 459527
rect 287713 459221 287747 459255
rect 296637 459493 296671 459527
rect 296637 459221 296671 459255
rect 306389 459493 306423 459527
rect 306389 459221 306423 459255
rect 315957 459493 315991 459527
rect 315957 459221 315991 459255
rect 331229 459289 331263 459323
rect 254961 459085 254995 459119
rect 332149 459289 332183 459323
rect 332149 459017 332183 459051
rect 334173 459289 334207 459323
rect 331229 458949 331263 458983
rect 334173 458881 334207 458915
rect 335369 459289 335403 459323
rect 249625 458813 249659 458847
rect 335369 458745 335403 458779
rect 337301 459289 337335 459323
rect 337301 458677 337335 458711
rect 338405 459289 338439 459323
rect 338405 458609 338439 458643
rect 340705 459289 340739 459323
rect 246497 458541 246531 458575
rect 243369 458473 243403 458507
rect 340705 458405 340739 458439
rect 341533 459289 341567 459323
rect 341533 458337 341567 458371
rect 240057 458269 240091 458303
rect 238033 458201 238067 458235
rect 317889 340153 317923 340187
rect 317889 338113 317923 338147
rect 326445 337501 326479 337535
rect 326261 337433 326295 337467
rect 331137 337433 331171 337467
rect 107485 336685 107519 336719
rect 100677 328389 100711 328423
rect 279525 336685 279559 336719
rect 331137 336685 331171 336719
rect 331229 337433 331263 337467
rect 331229 336685 331263 336719
rect 232145 335733 232179 335767
rect 232145 328457 232179 328491
rect 244473 334441 244507 334475
rect 244473 328457 244507 328491
rect 262781 333693 262815 333727
rect 107485 327097 107519 327131
rect 231133 328389 231167 328423
rect 100677 318801 100711 318835
rect 231133 318801 231167 318835
rect 254685 328389 254719 328423
rect 254685 318801 254719 318835
rect 257077 327029 257111 327063
rect 320281 335189 320315 335223
rect 279525 327097 279559 327131
rect 280629 328389 280663 328423
rect 262781 325669 262815 325703
rect 280629 318801 280663 318835
rect 281917 328389 281951 328423
rect 319453 328389 319487 328423
rect 295625 327029 295659 327063
rect 319453 325669 319487 325703
rect 344293 328389 344327 328423
rect 320281 325669 320315 325703
rect 341625 327029 341659 327063
rect 295625 322201 295659 322235
rect 335829 325601 335863 325635
rect 281917 318801 281951 318835
rect 257077 317441 257111 317475
rect 282653 318665 282687 318699
rect 107485 317373 107519 317407
rect 100677 309077 100711 309111
rect 244381 317373 244415 317407
rect 260389 317373 260423 317407
rect 244381 311457 244415 311491
rect 258825 315945 258859 315979
rect 107485 307785 107519 307819
rect 238033 309077 238067 309111
rect 100677 299489 100711 299523
rect 238033 299489 238067 299523
rect 257077 302889 257111 302923
rect 231225 299421 231259 299455
rect 107485 298061 107519 298095
rect 100677 289765 100711 289799
rect 240701 299421 240735 299455
rect 231225 289833 231259 289867
rect 232421 298061 232455 298095
rect 107485 288405 107519 288439
rect 240701 289833 240735 289867
rect 245025 298061 245059 298095
rect 232421 288405 232455 288439
rect 238033 289765 238067 289799
rect 100677 280177 100711 280211
rect 238033 280177 238067 280211
rect 231225 280109 231259 280143
rect 231225 270521 231259 270555
rect 240701 280109 240735 280143
rect 260389 307785 260423 307819
rect 261585 317373 261619 317407
rect 265817 317373 265851 317407
rect 344293 318801 344327 318835
rect 341625 317441 341659 317475
rect 335829 316013 335863 316047
rect 339969 317373 340003 317407
rect 319453 315945 319487 315979
rect 282653 309145 282687 309179
rect 293417 309145 293451 309179
rect 265817 307853 265851 307887
rect 261585 299489 261619 299523
rect 264529 307717 264563 307751
rect 258825 298129 258859 298163
rect 260297 299421 260331 299455
rect 257077 294457 257111 294491
rect 264529 298129 264563 298163
rect 265817 307717 265851 307751
rect 293417 306357 293451 306391
rect 316877 307717 316911 307751
rect 265817 298129 265851 298163
rect 319453 306357 319487 306391
rect 320281 315945 320315 315979
rect 339969 307785 340003 307819
rect 320281 306357 320315 306391
rect 316877 298129 316911 298163
rect 260297 289833 260331 289867
rect 319637 298061 319671 298095
rect 246405 288337 246439 288371
rect 245025 278749 245059 278783
rect 246037 280109 246071 280143
rect 240701 270521 240735 270555
rect 265817 288337 265851 288371
rect 258733 286977 258767 287011
rect 246405 278749 246439 278783
rect 257169 280109 257203 280143
rect 257169 278749 257203 278783
rect 321109 298061 321143 298095
rect 339969 298061 340003 298095
rect 321109 288473 321143 288507
rect 333161 289969 333195 290003
rect 333161 288405 333195 288439
rect 319637 287045 319671 287079
rect 339969 282829 340003 282863
rect 265817 278817 265851 278851
rect 258733 277389 258767 277423
rect 264529 278681 264563 278715
rect 246037 270521 246071 270555
rect 260297 273241 260331 273275
rect 100677 270453 100711 270487
rect 100677 260865 100711 260899
rect 238033 270453 238067 270487
rect 264529 269093 264563 269127
rect 265817 278681 265851 278715
rect 265817 269093 265851 269127
rect 260297 265285 260331 265319
rect 238033 260865 238067 260899
rect 322305 263585 322339 263619
rect 231225 260797 231259 260831
rect 322305 259437 322339 259471
rect 341625 260797 341659 260831
rect 232145 258009 232179 258043
rect 232145 253861 232179 253895
rect 232421 258009 232455 258043
rect 232421 253181 232455 253215
rect 244381 258009 244415 258043
rect 231225 251209 231259 251243
rect 100677 251141 100711 251175
rect 319637 258009 319671 258043
rect 299029 256649 299063 256683
rect 256985 251209 257019 251243
rect 256985 249781 257019 249815
rect 258825 249713 258859 249747
rect 244381 241553 244415 241587
rect 246313 248353 246347 248387
rect 100677 241485 100711 241519
rect 232697 240057 232731 240091
rect 299029 247061 299063 247095
rect 258825 240193 258859 240227
rect 300317 246993 300351 247027
rect 246313 238765 246347 238799
rect 232697 235297 232731 235331
rect 261585 238697 261619 238731
rect 232053 234617 232087 234651
rect 300317 237405 300351 237439
rect 301789 246993 301823 247027
rect 335737 258009 335771 258043
rect 334541 256649 334575 256683
rect 326261 254065 326295 254099
rect 334541 251073 334575 251107
rect 341625 251209 341659 251243
rect 335737 250937 335771 250971
rect 326261 249781 326295 249815
rect 319637 240125 319671 240159
rect 301789 237405 301823 237439
rect 261585 234549 261619 234583
rect 299029 237337 299063 237371
rect 232053 230469 232087 230503
rect 260389 229041 260423 229075
rect 232053 224961 232087 224995
rect 299029 227749 299063 227783
rect 301789 235909 301823 235943
rect 300317 227681 300351 227715
rect 260389 224213 260423 224247
rect 299029 227613 299063 227647
rect 232053 222173 232087 222207
rect 260389 219385 260423 219419
rect 246405 217413 246439 217447
rect 261585 219385 261619 219419
rect 299029 218025 299063 218059
rect 330401 235909 330435 235943
rect 330401 230061 330435 230095
rect 340061 229041 340095 229075
rect 301789 226321 301823 226355
rect 333069 227681 333103 227715
rect 300317 218025 300351 218059
rect 319637 219385 319671 219419
rect 261585 215237 261619 215271
rect 301789 216597 301823 216631
rect 260389 214489 260423 214523
rect 246405 209797 246439 209831
rect 300317 208301 300351 208335
rect 244473 202861 244507 202895
rect 244473 201501 244507 201535
rect 319637 209797 319671 209831
rect 321109 219385 321143 219419
rect 321109 209797 321143 209831
rect 322121 219317 322155 219351
rect 340061 220745 340095 220779
rect 333069 218025 333103 218059
rect 334633 216597 334667 216631
rect 322121 209797 322155 209831
rect 326261 215373 326295 215407
rect 301789 207009 301823 207043
rect 329021 215237 329055 215271
rect 340061 211089 340095 211123
rect 334633 207009 334667 207043
rect 335829 209729 335863 209763
rect 329021 205649 329055 205683
rect 326261 200141 326295 200175
rect 330585 205581 330619 205615
rect 300317 198713 300351 198747
rect 319637 200073 319671 200107
rect 299029 198645 299063 198679
rect 244933 195245 244967 195279
rect 244381 189465 244415 189499
rect 232329 182121 232363 182155
rect 244933 183549 244967 183583
rect 260205 191777 260239 191811
rect 260205 183481 260239 183515
rect 261493 190417 261527 190451
rect 244381 173893 244415 173927
rect 260297 182121 260331 182155
rect 261493 182121 261527 182155
rect 263057 190417 263091 190451
rect 299029 189057 299063 189091
rect 301789 197149 301823 197183
rect 263057 180829 263091 180863
rect 300317 188989 300351 189023
rect 260297 173825 260331 173859
rect 264529 180761 264563 180795
rect 232329 172533 232363 172567
rect 264529 171105 264563 171139
rect 265817 180761 265851 180795
rect 265817 171105 265851 171139
rect 293141 180761 293175 180795
rect 319637 190485 319671 190519
rect 321109 200073 321143 200107
rect 321109 190485 321143 190519
rect 322213 200073 322247 200107
rect 322213 190485 322247 190519
rect 329021 197285 329055 197319
rect 301789 187697 301823 187731
rect 329021 187697 329055 187731
rect 340061 204901 340095 204935
rect 335829 203541 335863 203575
rect 330585 187697 330619 187731
rect 334633 197285 334667 197319
rect 334633 187697 334667 187731
rect 335829 190417 335863 190451
rect 333161 183889 333195 183923
rect 333161 182053 333195 182087
rect 334541 180829 334575 180863
rect 335829 180829 335863 180863
rect 300317 179401 300351 179435
rect 319637 180761 319671 180795
rect 293141 171105 293175 171139
rect 301789 177973 301823 178007
rect 299029 169677 299063 169711
rect 107485 162809 107519 162843
rect 107485 153221 107519 153255
rect 232605 161381 232639 161415
rect 232053 153153 232087 153187
rect 232605 153153 232639 153187
rect 253029 161381 253063 161415
rect 253029 151793 253063 151827
rect 257077 161381 257111 161415
rect 293325 161381 293359 161415
rect 257077 151793 257111 151827
rect 260297 158661 260331 158695
rect 253029 151657 253063 151691
rect 232053 143565 232087 143599
rect 246405 143565 246439 143599
rect 107485 143497 107519 143531
rect 240701 143497 240735 143531
rect 232053 142069 232087 142103
rect 231225 137989 231259 138023
rect 231225 135337 231259 135371
rect 107485 133909 107519 133943
rect 232053 132481 232087 132515
rect 232421 136425 232455 136459
rect 107485 124117 107519 124151
rect 100677 115889 100711 115923
rect 246037 143497 246071 143531
rect 240701 133909 240735 133943
rect 244933 140709 244967 140743
rect 299029 160089 299063 160123
rect 300317 169677 300351 169711
rect 319637 171105 319671 171139
rect 321109 180761 321143 180795
rect 334541 179469 334575 179503
rect 321109 171105 321143 171139
rect 334541 179333 334575 179367
rect 334541 171037 334575 171071
rect 331781 169813 331815 169847
rect 301789 168385 301823 168419
rect 326353 169677 326387 169711
rect 300317 160089 300351 160123
rect 319637 161381 319671 161415
rect 293325 151793 293359 151827
rect 319637 151793 319671 151827
rect 321109 161381 321143 161415
rect 331781 168385 331815 168419
rect 326353 161313 326387 161347
rect 321109 151793 321143 151827
rect 260297 149073 260331 149107
rect 264529 151725 264563 151759
rect 253029 142205 253063 142239
rect 258825 143497 258859 143531
rect 246405 142137 246439 142171
rect 246037 133297 246071 133331
rect 246405 141865 246439 141899
rect 244933 131189 244967 131223
rect 253213 140709 253247 140743
rect 331781 151725 331815 151759
rect 264529 142137 264563 142171
rect 296085 150365 296119 150399
rect 293325 142069 293359 142103
rect 258825 138601 258859 138635
rect 260205 139349 260239 139383
rect 253213 131121 253247 131155
rect 330493 150365 330527 150399
rect 301513 150229 301547 150263
rect 301513 147645 301547 147679
rect 314393 143497 314427 143531
rect 296085 140777 296119 140811
rect 301881 141049 301915 141083
rect 293325 132481 293359 132515
rect 299029 140709 299063 140743
rect 260205 129761 260239 129795
rect 261493 131053 261527 131087
rect 246405 124185 246439 124219
rect 231225 118677 231259 118711
rect 232421 118677 232455 118711
rect 244381 122757 244415 122791
rect 231225 116025 231259 116059
rect 107485 114529 107519 114563
rect 231225 115889 231259 115923
rect 100677 106301 100711 106335
rect 253121 122757 253155 122791
rect 244381 113169 244415 113203
rect 245025 121397 245059 121431
rect 245025 113101 245059 113135
rect 244381 113033 244415 113067
rect 231225 106301 231259 106335
rect 232329 106981 232363 107015
rect 107485 104805 107519 104839
rect 100677 96577 100711 96611
rect 232145 102085 232179 102119
rect 231225 99365 231259 99399
rect 231225 96713 231259 96747
rect 107485 95217 107519 95251
rect 253121 108341 253155 108375
rect 254685 122757 254719 122791
rect 257169 122757 257203 122791
rect 300317 140709 300351 140743
rect 301881 140641 301915 140675
rect 314393 138465 314427 138499
rect 319637 142069 319671 142103
rect 300317 130713 300351 130747
rect 301789 134521 301823 134555
rect 299029 129829 299063 129863
rect 299029 129693 299063 129727
rect 261493 122689 261527 122723
rect 264621 122757 264655 122791
rect 261493 121261 261527 121295
rect 257169 113169 257203 113203
rect 258917 115889 258951 115923
rect 258917 106301 258951 106335
rect 260389 115889 260423 115923
rect 261493 111809 261527 111843
rect 263057 117997 263091 118031
rect 260389 106301 260423 106335
rect 254685 104873 254719 104907
rect 264621 113169 264655 113203
rect 265817 122757 265851 122791
rect 331781 142137 331815 142171
rect 334541 151725 334575 151759
rect 334541 142137 334575 142171
rect 330493 140777 330527 140811
rect 319637 132481 319671 132515
rect 329021 140709 329055 140743
rect 329021 131121 329055 131155
rect 331781 140709 331815 140743
rect 331781 131121 331815 131155
rect 335921 140709 335955 140743
rect 335921 131121 335955 131155
rect 340061 133841 340095 133875
rect 334449 131053 334483 131087
rect 301789 121465 301823 121499
rect 317153 124117 317187 124151
rect 299029 120173 299063 120207
rect 265817 113169 265851 113203
rect 298937 120037 298971 120071
rect 263057 104873 263091 104907
rect 294797 113101 294831 113135
rect 244381 103581 244415 103615
rect 294797 103513 294831 103547
rect 297465 106913 297499 106947
rect 253213 103445 253247 103479
rect 246313 99433 246347 99467
rect 246313 95149 246347 95183
rect 258917 103445 258951 103479
rect 253213 95149 253247 95183
rect 257077 95149 257111 95183
rect 232329 93857 232363 93891
rect 232145 92497 232179 92531
rect 100677 86989 100711 87023
rect 232329 89709 232363 89743
rect 107485 85493 107519 85527
rect 100677 77197 100711 77231
rect 107485 75905 107519 75939
rect 253029 85629 253063 85663
rect 263057 103445 263091 103479
rect 258917 93857 258951 93891
rect 261585 99773 261619 99807
rect 257077 85561 257111 85595
rect 263057 93857 263091 93891
rect 264437 103445 264471 103479
rect 265725 103445 265759 103479
rect 265725 95149 265759 95183
rect 293325 103445 293359 103479
rect 264437 93857 264471 93891
rect 298937 102153 298971 102187
rect 300225 120037 300259 120071
rect 300225 102153 300259 102187
rect 301697 120037 301731 120071
rect 317153 117521 317187 117555
rect 317337 124117 317371 124151
rect 317337 115549 317371 115583
rect 319637 122621 319671 122655
rect 316969 114461 317003 114495
rect 317153 114461 317187 114495
rect 317337 114461 317371 114495
rect 317153 107593 317187 107627
rect 317245 114393 317279 114427
rect 340061 124185 340095 124219
rect 334449 121465 334483 121499
rect 319637 113169 319671 113203
rect 331781 121397 331815 121431
rect 317337 109701 317371 109735
rect 326169 113101 326203 113135
rect 317245 106097 317279 106131
rect 316969 104873 317003 104907
rect 321109 106029 321143 106063
rect 301697 102153 301731 102187
rect 319637 103445 319671 103479
rect 297465 100725 297499 100759
rect 293325 93857 293359 93891
rect 319637 93857 319671 93891
rect 339969 115481 340003 115515
rect 331781 111809 331815 111843
rect 335829 113101 335863 113135
rect 326169 103513 326203 103547
rect 334541 111741 334575 111775
rect 321109 93857 321143 93891
rect 322305 103445 322339 103479
rect 339969 108953 340003 108987
rect 335829 103581 335863 103615
rect 334541 102221 334575 102255
rect 335921 103445 335955 103479
rect 322305 93857 322339 93891
rect 328929 102085 328963 102119
rect 328929 92497 328963 92531
rect 334541 102085 334575 102119
rect 335921 93857 335955 93891
rect 340061 95149 340095 95183
rect 334541 92497 334575 92531
rect 296637 89029 296671 89063
rect 296637 86853 296671 86887
rect 340061 85561 340095 85595
rect 261585 85493 261619 85527
rect 253029 84201 253063 84235
rect 320833 84269 320867 84303
rect 244473 84133 244507 84167
rect 261677 84133 261711 84167
rect 244473 77197 244507 77231
rect 246037 77333 246071 77367
rect 232329 75905 232363 75939
rect 246037 74545 246071 74579
rect 254777 75837 254811 75871
rect 253213 73117 253247 73151
rect 100677 67609 100711 67643
rect 232145 73049 232179 73083
rect 107485 66181 107519 66215
rect 100677 57885 100711 57919
rect 107485 56593 107519 56627
rect 100677 48297 100711 48331
rect 231317 55165 231351 55199
rect 107485 46869 107519 46903
rect 100677 38573 100711 38607
rect 264529 84133 264563 84167
rect 261677 74613 261711 74647
rect 263057 82977 263091 83011
rect 254777 69649 254811 69683
rect 264529 74545 264563 74579
rect 293325 84133 293359 84167
rect 293325 74545 293359 74579
rect 294797 84133 294831 84167
rect 319637 84133 319671 84167
rect 294797 74545 294831 74579
rect 314209 77197 314243 77231
rect 263057 67609 263091 67643
rect 314209 67609 314243 67643
rect 318165 77197 318199 77231
rect 320833 82909 320867 82943
rect 319637 74545 319671 74579
rect 320833 82773 320867 82807
rect 320833 73185 320867 73219
rect 329021 82773 329055 82807
rect 329021 71757 329055 71791
rect 318165 67609 318199 67643
rect 345397 67541 345431 67575
rect 314209 66181 314243 66215
rect 253213 63529 253247 63563
rect 264529 64821 264563 64855
rect 254777 63461 254811 63495
rect 246497 57885 246531 57919
rect 240609 56525 240643 56559
rect 240609 47005 240643 47039
rect 244473 56525 244507 56559
rect 232145 46937 232179 46971
rect 254777 53805 254811 53839
rect 261585 55981 261619 56015
rect 246497 48297 246531 48331
rect 244473 46937 244507 46971
rect 261585 46937 261619 46971
rect 265817 64821 265851 64855
rect 265817 55301 265851 55335
rect 293325 64821 293359 64855
rect 264529 46937 264563 46971
rect 265817 55165 265851 55199
rect 231317 45577 231351 45611
rect 240701 46869 240735 46903
rect 107485 37281 107519 37315
rect 232329 40681 232363 40715
rect 100677 28985 100711 29019
rect 232329 27625 232363 27659
rect 232789 40681 232823 40715
rect 293325 46937 293359 46971
rect 294797 64821 294831 64855
rect 294797 46937 294831 46971
rect 296085 59993 296119 60027
rect 314209 56593 314243 56627
rect 319637 64821 319671 64855
rect 296085 46937 296119 46971
rect 299029 55165 299063 55199
rect 265817 45577 265851 45611
rect 299029 45577 299063 45611
rect 300317 55165 300351 55199
rect 300317 45577 300351 45611
rect 301789 55165 301823 55199
rect 322305 64821 322339 64855
rect 319637 46937 319671 46971
rect 321017 63461 321051 63495
rect 301789 45577 301823 45611
rect 314209 46869 314243 46903
rect 252937 45509 252971 45543
rect 244381 41429 244415 41463
rect 252937 40681 252971 40715
rect 257169 45509 257203 45543
rect 244381 38573 244415 38607
rect 240701 37349 240735 37383
rect 232789 27625 232823 27659
rect 252937 35853 252971 35887
rect 107485 27557 107519 27591
rect 244473 27557 244507 27591
rect 264437 45509 264471 45543
rect 261585 42109 261619 42143
rect 261585 35921 261619 35955
rect 264437 35921 264471 35955
rect 265725 37349 265759 37383
rect 322305 55301 322339 55335
rect 331781 63461 331815 63495
rect 331781 53805 331815 53839
rect 334541 61421 334575 61455
rect 345397 57953 345431 57987
rect 334541 46937 334575 46971
rect 321017 45577 321051 45611
rect 314209 37281 314243 37315
rect 319637 45509 319671 45543
rect 265725 35921 265759 35955
rect 322305 45509 322339 45543
rect 319637 35921 319671 35955
rect 321017 40681 321051 40715
rect 322305 40681 322339 40715
rect 326353 44081 326387 44115
rect 257169 27625 257203 27659
rect 299029 35853 299063 35887
rect 252937 26265 252971 26299
rect 299029 26265 299063 26299
rect 300317 35853 300351 35887
rect 300317 26265 300351 26299
rect 301789 35853 301823 35887
rect 321017 31705 321051 31739
rect 326353 27625 326387 27659
rect 301789 26265 301823 26299
rect 314209 27557 314243 27591
rect 300685 23409 300719 23443
rect 244473 17969 244507 18003
rect 297557 23341 297591 23375
rect 278421 17153 278455 17187
rect 278237 17085 278271 17119
rect 268761 16677 268795 16711
rect 231133 16541 231167 16575
rect 231409 16541 231443 16575
rect 268945 16677 268979 16711
rect 268761 13073 268795 13107
rect 268853 16609 268887 16643
rect 268945 13141 268979 13175
rect 269037 16609 269071 16643
rect 269037 13073 269071 13107
rect 278329 17085 278363 17119
rect 278329 12801 278363 12835
rect 278237 12733 278271 12767
rect 268853 12529 268887 12563
rect 107485 9673 107519 9707
rect 278605 17153 278639 17187
rect 90925 9605 90959 9639
rect 58725 4097 58759 4131
rect 55229 3825 55263 3859
rect 55229 3689 55263 3723
rect 34621 3621 34655 3655
rect 34621 3349 34655 3383
rect 55229 3553 55263 3587
rect 55229 3281 55263 3315
rect 55321 3213 55355 3247
rect 58725 3349 58759 3383
rect 64797 3825 64831 3859
rect 55413 3145 55447 3179
rect 64797 3689 64831 3723
rect 64889 3621 64923 3655
rect 64797 3553 64831 3587
rect 64705 3281 64739 3315
rect 64613 3213 64647 3247
rect 64521 3145 64555 3179
rect 64889 3145 64923 3179
rect 74457 3621 74491 3655
rect 74457 3145 74491 3179
rect 84209 3621 84243 3655
rect 84209 3009 84243 3043
rect 100493 9605 100527 9639
rect 99297 3621 99331 3655
rect 99297 2941 99331 2975
rect 90925 561 90959 595
rect 108773 9605 108807 9639
rect 278421 9605 278455 9639
rect 278513 17085 278547 17119
rect 101505 3621 101539 3655
rect 101505 2805 101539 2839
rect 100493 561 100527 595
rect 278697 17085 278731 17119
rect 301789 18241 301823 18275
rect 301789 14365 301823 14399
rect 301881 18173 301915 18207
rect 304641 18037 304675 18071
rect 302065 17289 302099 17323
rect 301973 17221 302007 17255
rect 301973 15181 302007 15215
rect 302157 17221 302191 17255
rect 302157 15181 302191 15215
rect 304641 15181 304675 15215
rect 304917 17969 304951 18003
rect 314209 17969 314243 18003
rect 329113 17969 329147 18003
rect 304917 15181 304951 15215
rect 307217 15181 307251 15215
rect 329113 15181 329147 15215
rect 302065 15113 302099 15147
rect 301881 14297 301915 14331
rect 300685 14025 300719 14059
rect 297557 13957 297591 13991
rect 278697 13073 278731 13107
rect 278605 12053 278639 12087
rect 307217 11373 307251 11407
rect 278513 9537 278547 9571
rect 345397 11033 345431 11067
rect 323133 9129 323167 9163
rect 322673 9061 322707 9095
rect 323041 9061 323075 9095
rect 322765 8993 322799 9027
rect 324513 8993 324547 9027
rect 324053 8925 324087 8959
rect 345397 8313 345431 8347
rect 252937 8245 252971 8279
rect 250269 5525 250303 5559
rect 135269 4709 135303 4743
rect 135453 4709 135487 4743
rect 154589 4709 154623 4743
rect 154773 4709 154807 4743
rect 135177 4641 135211 4675
rect 125609 4573 125643 4607
rect 125609 4437 125643 4471
rect 135361 4641 135395 4675
rect 154497 4641 154531 4675
rect 135361 4505 135395 4539
rect 144929 4505 144963 4539
rect 135177 4437 135211 4471
rect 144929 4369 144963 4403
rect 154497 4369 154531 4403
rect 154589 4573 154623 4607
rect 238769 4573 238803 4607
rect 239689 4573 239723 4607
rect 246681 4573 246715 4607
rect 154589 4369 154623 4403
rect 164157 4505 164191 4539
rect 239045 4505 239079 4539
rect 239413 4505 239447 4539
rect 246681 4437 246715 4471
rect 280077 6341 280111 6375
rect 252937 5389 252971 5423
rect 267289 5525 267323 5559
rect 268393 5525 268427 5559
rect 267289 5321 267323 5355
rect 268301 5321 268335 5355
rect 268393 5321 268427 5355
rect 268301 4913 268335 4947
rect 270693 5049 270727 5083
rect 267381 4845 267415 4879
rect 264989 4777 265023 4811
rect 250269 4437 250303 4471
rect 263425 4505 263459 4539
rect 164157 4369 164191 4403
rect 263425 4369 263459 4403
rect 264989 4369 265023 4403
rect 176577 4301 176611 4335
rect 128277 4165 128311 4199
rect 117329 3621 117363 3655
rect 119353 3621 119387 3655
rect 124229 3621 124263 3655
rect 128277 3621 128311 3655
rect 128369 4165 128403 4199
rect 128369 3621 128403 3655
rect 147597 4165 147631 4199
rect 147597 3621 147631 3655
rect 157257 4165 157291 4199
rect 176485 4165 176519 4199
rect 157257 3621 157291 3655
rect 168665 3553 168699 3587
rect 168757 3825 168791 3859
rect 168849 3825 168883 3859
rect 171701 3825 171735 3859
rect 171793 3825 171827 3859
rect 171793 3621 171827 3655
rect 168757 3553 168791 3587
rect 171793 3349 171827 3383
rect 171885 3349 171919 3383
rect 171977 3689 172011 3723
rect 215125 4301 215159 4335
rect 180717 4165 180751 4199
rect 180625 3825 180659 3859
rect 176577 3621 176611 3655
rect 180533 3689 180567 3723
rect 176485 3349 176519 3383
rect 180625 3553 180659 3587
rect 180809 4165 180843 4199
rect 180809 3621 180843 3655
rect 190377 4165 190411 4199
rect 190377 3621 190411 3655
rect 200129 4165 200163 4199
rect 205741 4165 205775 4199
rect 205741 3689 205775 3723
rect 215033 4165 215067 4199
rect 200129 3621 200163 3655
rect 180717 3553 180751 3587
rect 208041 3553 208075 3587
rect 180717 3349 180751 3383
rect 208133 3553 208167 3587
rect 215493 4301 215527 4335
rect 215217 4233 215251 4267
rect 215217 3825 215251 3859
rect 215309 4233 215343 4267
rect 215309 3825 215343 3859
rect 215401 4165 215435 4199
rect 215401 3689 215435 3723
rect 215125 3621 215159 3655
rect 208133 3349 208167 3383
rect 208225 3349 208259 3383
rect 215033 3349 215067 3383
rect 239505 4301 239539 4335
rect 264805 4301 264839 4335
rect 265081 4301 265115 4335
rect 267381 4301 267415 4335
rect 268393 4709 268427 4743
rect 270693 4709 270727 4743
rect 270785 4709 270819 4743
rect 268393 4233 268427 4267
rect 220185 4165 220219 4199
rect 224877 4165 224911 4199
rect 239229 4165 239263 4199
rect 270785 4165 270819 4199
rect 220185 3689 220219 3723
rect 220277 3689 220311 3723
rect 220093 3553 220127 3587
rect 215493 3349 215527 3383
rect 220001 3349 220035 3383
rect 220093 3349 220127 3383
rect 263609 3825 263643 3859
rect 224877 3553 224911 3587
rect 270509 3621 270543 3655
rect 263701 3553 263735 3587
rect 266001 3553 266035 3587
rect 266093 3553 266127 3587
rect 266093 3349 266127 3383
rect 266185 3349 266219 3383
rect 267749 3349 267783 3383
rect 270509 3349 270543 3383
rect 277317 3349 277351 3383
rect 277961 3349 277995 3383
rect 278053 3553 278087 3587
rect 278145 3553 278179 3587
rect 278053 3349 278087 3383
rect 119353 2941 119387 2975
rect 124137 2941 124171 2975
rect 124229 2941 124263 2975
rect 117053 2805 117087 2839
rect 124229 2737 124263 2771
rect 267749 2737 267783 2771
rect 277317 2737 277351 2771
rect 108773 561 108807 595
rect 292497 4301 292531 4335
rect 282745 4233 282779 4267
rect 292405 4233 292439 4267
rect 282745 3825 282779 3859
rect 282837 3825 282871 3859
rect 282745 3553 282779 3587
rect 285321 3553 285355 3587
rect 285413 3553 285447 3587
rect 285413 3349 285447 3383
rect 285505 3349 285539 3383
rect 292497 3825 292531 3859
rect 292589 4301 292623 4335
rect 292589 3825 292623 3859
rect 292681 4233 292715 4267
rect 292405 3349 292439 3383
rect 326537 4165 326571 4199
rect 303997 3825 304031 3859
rect 304089 3825 304123 3859
rect 306941 3825 306975 3859
rect 307033 3825 307067 3859
rect 303813 3689 303847 3723
rect 303905 3689 303939 3723
rect 297373 3553 297407 3587
rect 292681 3349 292715 3383
rect 297281 3349 297315 3383
rect 297373 3349 297407 3383
rect 297465 3553 297499 3587
rect 303905 3553 303939 3587
rect 303997 3553 304031 3587
rect 306849 3689 306883 3723
rect 306941 3689 306975 3723
rect 307033 3621 307067 3655
rect 316693 3825 316727 3859
rect 316785 3825 316819 3859
rect 313749 3689 313783 3723
rect 307125 3621 307159 3655
rect 313657 3621 313691 3655
rect 306941 3349 306975 3383
rect 307033 3349 307067 3383
rect 313657 3349 313691 3383
rect 324973 3689 325007 3723
rect 317061 3621 317095 3655
rect 316785 3553 316819 3587
rect 326261 3621 326295 3655
rect 326629 3621 326663 3655
rect 324973 3485 325007 3519
rect 313749 3349 313783 3383
rect 326629 3349 326663 3383
rect 280077 561 280111 595
<< metal1 >>
rect 170306 700952 170312 701004
rect 170364 700992 170370 701004
rect 293218 700992 293224 701004
rect 170364 700964 293224 700992
rect 170364 700952 170370 700964
rect 293218 700952 293224 700964
rect 293276 700952 293282 701004
rect 286962 700884 286968 700936
rect 287020 700924 287026 700936
rect 413646 700924 413652 700936
rect 287020 700896 413652 700924
rect 287020 700884 287026 700896
rect 413646 700884 413652 700896
rect 413704 700884 413710 700936
rect 284202 700816 284208 700868
rect 284260 700856 284266 700868
rect 429838 700856 429844 700868
rect 284260 700828 429844 700856
rect 284260 700816 284266 700828
rect 429838 700816 429844 700828
rect 429896 700816 429902 700868
rect 137830 700748 137836 700800
rect 137888 700788 137894 700800
rect 294598 700788 294604 700800
rect 137888 700760 294604 700788
rect 137888 700748 137894 700760
rect 294598 700748 294604 700760
rect 294656 700748 294662 700800
rect 282822 700680 282828 700732
rect 282880 700720 282886 700732
rect 462314 700720 462320 700732
rect 282880 700692 462320 700720
rect 282880 700680 282886 700692
rect 462314 700680 462320 700692
rect 462372 700680 462378 700732
rect 105446 700612 105452 700664
rect 105504 700652 105510 700664
rect 295978 700652 295984 700664
rect 105504 700624 295984 700652
rect 105504 700612 105510 700624
rect 295978 700612 295984 700624
rect 296036 700612 296042 700664
rect 284110 700544 284116 700596
rect 284168 700584 284174 700596
rect 478506 700584 478512 700596
rect 284168 700556 478512 700584
rect 284168 700544 284174 700556
rect 478506 700544 478512 700556
rect 478564 700544 478570 700596
rect 72970 700476 72976 700528
rect 73028 700516 73034 700528
rect 297358 700516 297364 700528
rect 73028 700488 297364 700516
rect 73028 700476 73034 700488
rect 297358 700476 297364 700488
rect 297416 700476 297422 700528
rect 299474 700476 299480 700528
rect 299532 700516 299538 700528
rect 300118 700516 300124 700528
rect 299532 700488 300124 700516
rect 299532 700476 299538 700488
rect 300118 700476 300124 700488
rect 300176 700476 300182 700528
rect 280062 700408 280068 700460
rect 280120 700448 280126 700460
rect 527174 700448 527180 700460
rect 280120 700420 527180 700448
rect 280120 700408 280126 700420
rect 527174 700408 527180 700420
rect 527232 700408 527238 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 300118 700380 300124 700392
rect 40552 700352 300124 700380
rect 40552 700340 40558 700352
rect 300118 700340 300124 700352
rect 300176 700340 300182 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 301498 700312 301504 700324
rect 8168 700284 301504 700312
rect 8168 700272 8174 700284
rect 301498 700272 301504 700284
rect 301556 700272 301562 700324
rect 285582 700204 285588 700256
rect 285640 700244 285646 700256
rect 397454 700244 397460 700256
rect 285640 700216 397460 700244
rect 285640 700204 285646 700216
rect 397454 700204 397460 700216
rect 397512 700204 397518 700256
rect 202782 700136 202788 700188
rect 202840 700176 202846 700188
rect 291838 700176 291844 700188
rect 202840 700148 291844 700176
rect 202840 700136 202846 700148
rect 291838 700136 291844 700148
rect 291896 700136 291902 700188
rect 288342 700068 288348 700120
rect 288400 700108 288406 700120
rect 364978 700108 364984 700120
rect 288400 700080 364984 700108
rect 288400 700068 288406 700080
rect 364978 700068 364984 700080
rect 365036 700068 365042 700120
rect 289722 700000 289728 700052
rect 289780 700040 289786 700052
rect 348786 700040 348792 700052
rect 289780 700012 348792 700040
rect 289780 700000 289786 700012
rect 348786 700000 348792 700012
rect 348844 700000 348850 700052
rect 235166 699932 235172 699984
rect 235224 699972 235230 699984
rect 290458 699972 290464 699984
rect 235224 699944 290464 699972
rect 235224 699932 235230 699944
rect 290458 699932 290464 699944
rect 290516 699932 290522 699984
rect 291102 699932 291108 699984
rect 291160 699972 291166 699984
rect 299474 699972 299480 699984
rect 291160 699944 299480 699972
rect 291160 699932 291166 699944
rect 299474 699932 299480 699944
rect 299532 699932 299538 699984
rect 288250 699864 288256 699916
rect 288308 699904 288314 699916
rect 332502 699904 332508 699916
rect 288308 699876 332508 699904
rect 288308 699864 288314 699876
rect 332502 699864 332508 699876
rect 332560 699864 332566 699916
rect 283834 699796 283840 699848
rect 283892 699836 283898 699848
rect 291286 699836 291292 699848
rect 283892 699808 291292 699836
rect 283892 699796 283898 699808
rect 291286 699796 291292 699808
rect 291344 699796 291350 699848
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 89162 699660 89168 699712
rect 89220 699700 89226 699712
rect 89622 699700 89628 699712
rect 89220 699672 89628 699700
rect 89220 699660 89226 699672
rect 89622 699660 89628 699672
rect 89680 699660 89686 699712
rect 542722 698232 542728 698284
rect 542780 698272 542786 698284
rect 543550 698272 543556 698284
rect 542780 698244 543556 698272
rect 542780 698232 542786 698244
rect 543550 698232 543556 698244
rect 543608 698232 543614 698284
rect 275922 696940 275928 696992
rect 275980 696980 275986 696992
rect 580166 696980 580172 696992
rect 275980 696952 580172 696980
rect 275980 696940 275986 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 154114 695512 154120 695564
rect 154172 695552 154178 695564
rect 154206 695552 154212 695564
rect 154172 695524 154212 695552
rect 154172 695512 154178 695524
rect 154206 695512 154212 695524
rect 154264 695512 154270 695564
rect 218974 694152 218980 694204
rect 219032 694192 219038 694204
rect 219158 694192 219164 694204
rect 219032 694164 219164 694192
rect 219032 694152 219038 694164
rect 219158 694152 219164 694164
rect 219216 694152 219222 694204
rect 219158 688684 219164 688696
rect 219084 688656 219164 688684
rect 219084 688628 219112 688656
rect 219158 688644 219164 688656
rect 219216 688644 219222 688696
rect 542722 688644 542728 688696
rect 542780 688644 542786 688696
rect 154206 688576 154212 688628
rect 154264 688616 154270 688628
rect 154390 688616 154396 688628
rect 154264 688588 154396 688616
rect 154264 688576 154270 688588
rect 154390 688576 154396 688588
rect 154448 688576 154454 688628
rect 219066 688576 219072 688628
rect 219124 688576 219130 688628
rect 542538 688576 542544 688628
rect 542596 688616 542602 688628
rect 542740 688616 542768 688644
rect 542596 688588 542768 688616
rect 542596 688576 542602 688588
rect 559098 688576 559104 688628
rect 559156 688616 559162 688628
rect 559650 688616 559656 688628
rect 559156 688588 559656 688616
rect 559156 688576 559162 688588
rect 559650 688576 559656 688588
rect 559708 688576 559714 688628
rect 540992 685936 542860 685964
rect 277302 685856 277308 685908
rect 277360 685896 277366 685908
rect 540992 685896 541020 685936
rect 277360 685868 541020 685896
rect 542832 685896 542860 685936
rect 552584 685936 559788 685964
rect 552584 685896 552612 685936
rect 542832 685868 552612 685896
rect 559760 685896 559788 685936
rect 580166 685896 580172 685908
rect 559760 685868 580172 685896
rect 277360 685856 277366 685868
rect 580166 685856 580172 685868
rect 580224 685856 580230 685908
rect 154301 685831 154359 685837
rect 154301 685797 154313 685831
rect 154347 685828 154359 685831
rect 154390 685828 154396 685840
rect 154347 685800 154396 685828
rect 154347 685797 154359 685800
rect 154301 685791 154359 685797
rect 154390 685788 154396 685800
rect 154448 685788 154454 685840
rect 542446 684428 542452 684480
rect 542504 684468 542510 684480
rect 542725 684471 542783 684477
rect 542725 684468 542737 684471
rect 542504 684440 542737 684468
rect 542504 684428 542510 684440
rect 542725 684437 542737 684440
rect 542771 684437 542783 684471
rect 542725 684431 542783 684437
rect 559006 684428 559012 684480
rect 559064 684468 559070 684480
rect 559285 684471 559343 684477
rect 559285 684468 559297 684471
rect 559064 684440 559297 684468
rect 559064 684428 559070 684440
rect 559285 684437 559297 684440
rect 559331 684437 559343 684471
rect 559285 684431 559343 684437
rect 3510 681708 3516 681760
rect 3568 681748 3574 681760
rect 305086 681748 305092 681760
rect 3568 681720 305092 681748
rect 3568 681708 3574 681720
rect 305086 681708 305092 681720
rect 305144 681708 305150 681760
rect 154298 676240 154304 676252
rect 154259 676212 154304 676240
rect 154298 676200 154304 676212
rect 154356 676200 154362 676252
rect 218974 676172 218980 676184
rect 218935 676144 218980 676172
rect 218974 676132 218980 676144
rect 219032 676132 219038 676184
rect 494054 676172 494060 676184
rect 494015 676144 494060 676172
rect 494054 676132 494060 676144
rect 494112 676132 494118 676184
rect 154298 673480 154304 673532
rect 154356 673520 154362 673532
rect 154482 673520 154488 673532
rect 154356 673492 154488 673520
rect 154356 673480 154362 673492
rect 154482 673480 154488 673492
rect 154540 673480 154546 673532
rect 274542 673480 274548 673532
rect 274600 673520 274606 673532
rect 580166 673520 580172 673532
rect 274600 673492 580172 673520
rect 274600 673480 274606 673492
rect 580166 673480 580172 673492
rect 580224 673480 580230 673532
rect 3418 667904 3424 667956
rect 3476 667944 3482 667956
rect 305638 667944 305644 667956
rect 3476 667916 305644 667944
rect 3476 667904 3482 667916
rect 305638 667904 305644 667916
rect 305696 667904 305702 667956
rect 218977 666587 219035 666593
rect 218977 666553 218989 666587
rect 219023 666584 219035 666587
rect 219066 666584 219072 666596
rect 219023 666556 219072 666584
rect 219023 666553 219035 666556
rect 218977 666547 219035 666553
rect 219066 666544 219072 666556
rect 219124 666544 219130 666596
rect 494057 666587 494115 666593
rect 494057 666553 494069 666587
rect 494103 666584 494115 666587
rect 494146 666584 494152 666596
rect 494103 666556 494152 666584
rect 494103 666553 494115 666556
rect 494057 666547 494115 666553
rect 494146 666544 494152 666556
rect 494204 666544 494210 666596
rect 542725 666587 542783 666593
rect 542725 666553 542737 666587
rect 542771 666584 542783 666587
rect 542814 666584 542820 666596
rect 542771 666556 542820 666584
rect 542771 666553 542783 666556
rect 542725 666547 542783 666553
rect 542814 666544 542820 666556
rect 542872 666544 542878 666596
rect 559285 666587 559343 666593
rect 559285 666553 559297 666587
rect 559331 666584 559343 666587
rect 559374 666584 559380 666596
rect 559331 666556 559380 666584
rect 559331 666553 559343 666556
rect 559285 666547 559343 666553
rect 559374 666544 559380 666556
rect 559432 666544 559438 666596
rect 219158 659608 219164 659660
rect 219216 659648 219222 659660
rect 219342 659648 219348 659660
rect 219216 659620 219348 659648
rect 219216 659608 219222 659620
rect 219342 659608 219348 659620
rect 219400 659608 219406 659660
rect 219253 656863 219311 656869
rect 219253 656829 219265 656863
rect 219299 656860 219311 656863
rect 219342 656860 219348 656872
rect 219299 656832 219348 656860
rect 219299 656829 219311 656832
rect 219253 656823 219311 656829
rect 219342 656820 219348 656832
rect 219400 656820 219406 656872
rect 154298 654100 154304 654152
rect 154356 654140 154362 654152
rect 154482 654140 154488 654152
rect 154356 654112 154488 654140
rect 154356 654100 154362 654112
rect 154482 654100 154488 654112
rect 154540 654100 154546 654152
rect 494054 654100 494060 654152
rect 494112 654140 494118 654152
rect 494238 654140 494244 654152
rect 494112 654112 494244 654140
rect 494112 654100 494118 654112
rect 494238 654100 494244 654112
rect 494296 654100 494302 654152
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 306374 652780 306380 652792
rect 3108 652752 306380 652780
rect 3108 652740 3114 652752
rect 306374 652740 306380 652752
rect 306432 652740 306438 652792
rect 273162 650020 273168 650072
rect 273220 650060 273226 650072
rect 580166 650060 580172 650072
rect 273220 650032 580172 650060
rect 273220 650020 273226 650032
rect 580166 650020 580172 650032
rect 580224 650020 580230 650072
rect 219250 647272 219256 647284
rect 219211 647244 219256 647272
rect 219250 647232 219256 647244
rect 219308 647232 219314 647284
rect 542538 647232 542544 647284
rect 542596 647272 542602 647284
rect 542630 647272 542636 647284
rect 542596 647244 542636 647272
rect 542596 647232 542602 647244
rect 542630 647232 542636 647244
rect 542688 647232 542694 647284
rect 559098 647232 559104 647284
rect 559156 647272 559162 647284
rect 559190 647272 559196 647284
rect 559156 647244 559196 647272
rect 559156 647232 559162 647244
rect 559190 647232 559196 647244
rect 559248 647232 559254 647284
rect 219250 640404 219256 640416
rect 219084 640376 219256 640404
rect 219084 640280 219112 640376
rect 219250 640364 219256 640376
rect 219308 640364 219314 640416
rect 542538 640364 542544 640416
rect 542596 640404 542602 640416
rect 542630 640404 542636 640416
rect 542596 640376 542636 640404
rect 542596 640364 542602 640376
rect 542630 640364 542636 640376
rect 542688 640364 542694 640416
rect 559098 640364 559104 640416
rect 559156 640404 559162 640416
rect 559190 640404 559196 640416
rect 559156 640376 559196 640404
rect 559156 640364 559162 640376
rect 559190 640364 559196 640376
rect 559248 640364 559254 640416
rect 219066 640228 219072 640280
rect 219124 640228 219130 640280
rect 274450 638936 274456 638988
rect 274508 638976 274514 638988
rect 580166 638976 580172 638988
rect 274508 638948 580172 638976
rect 274508 638936 274514 638948
rect 580166 638936 580172 638948
rect 580224 638936 580230 638988
rect 219066 637508 219072 637560
rect 219124 637548 219130 637560
rect 219158 637548 219164 637560
rect 219124 637520 219164 637548
rect 219124 637508 219130 637520
rect 219158 637508 219164 637520
rect 219216 637508 219222 637560
rect 154298 634788 154304 634840
rect 154356 634828 154362 634840
rect 154482 634828 154488 634840
rect 154356 634800 154488 634828
rect 154356 634788 154362 634800
rect 154482 634788 154488 634800
rect 154540 634788 154546 634840
rect 494054 634788 494060 634840
rect 494112 634828 494118 634840
rect 494238 634828 494244 634840
rect 494112 634800 494244 634828
rect 494112 634788 494118 634800
rect 494238 634788 494244 634800
rect 494296 634788 494302 634840
rect 542446 630640 542452 630692
rect 542504 630680 542510 630692
rect 542630 630680 542636 630692
rect 542504 630652 542636 630680
rect 542504 630640 542510 630652
rect 542630 630640 542636 630652
rect 542688 630640 542694 630692
rect 559006 630640 559012 630692
rect 559064 630680 559070 630692
rect 559190 630680 559196 630692
rect 559064 630652 559196 630680
rect 559064 630640 559070 630652
rect 559190 630640 559196 630652
rect 559248 630640 559254 630692
rect 271782 626560 271788 626612
rect 271840 626600 271846 626612
rect 580166 626600 580172 626612
rect 271840 626572 580172 626600
rect 271840 626560 271846 626572
rect 580166 626560 580172 626572
rect 580224 626560 580230 626612
rect 219342 626532 219348 626544
rect 219303 626504 219348 626532
rect 219342 626492 219348 626504
rect 219400 626492 219406 626544
rect 3418 623772 3424 623824
rect 3476 623812 3482 623824
rect 309134 623812 309140 623824
rect 3476 623784 309140 623812
rect 3476 623772 3482 623784
rect 309134 623772 309140 623784
rect 309192 623772 309198 623824
rect 219342 616876 219348 616888
rect 219303 616848 219348 616876
rect 219342 616836 219348 616848
rect 219400 616836 219406 616888
rect 154298 615476 154304 615528
rect 154356 615516 154362 615528
rect 154482 615516 154488 615528
rect 154356 615488 154488 615516
rect 154356 615476 154362 615488
rect 154482 615476 154488 615488
rect 154540 615476 154546 615528
rect 494054 615476 494060 615528
rect 494112 615516 494118 615528
rect 494238 615516 494244 615528
rect 494112 615488 494244 615516
rect 494112 615476 494118 615488
rect 494238 615476 494244 615488
rect 494296 615476 494302 615528
rect 219069 611439 219127 611445
rect 219069 611405 219081 611439
rect 219115 611436 219127 611439
rect 219342 611436 219348 611448
rect 219115 611408 219348 611436
rect 219115 611405 219127 611408
rect 219069 611399 219127 611405
rect 219342 611396 219348 611408
rect 219400 611396 219406 611448
rect 542446 611328 542452 611380
rect 542504 611368 542510 611380
rect 542630 611368 542636 611380
rect 542504 611340 542636 611368
rect 542504 611328 542510 611340
rect 542630 611328 542636 611340
rect 542688 611328 542694 611380
rect 559006 611328 559012 611380
rect 559064 611368 559070 611380
rect 559190 611368 559196 611380
rect 559064 611340 559196 611368
rect 559064 611328 559070 611340
rect 559190 611328 559196 611340
rect 559248 611328 559254 611380
rect 3418 609968 3424 610020
rect 3476 610008 3482 610020
rect 308398 610008 308404 610020
rect 3476 609980 308404 610008
rect 3476 609968 3482 609980
rect 308398 609968 308404 609980
rect 308456 609968 308462 610020
rect 219066 608716 219072 608728
rect 219027 608688 219072 608716
rect 219066 608676 219072 608688
rect 219124 608676 219130 608728
rect 219066 608540 219072 608592
rect 219124 608580 219130 608592
rect 219253 608583 219311 608589
rect 219253 608580 219265 608583
rect 219124 608552 219265 608580
rect 219124 608540 219130 608552
rect 219253 608549 219265 608552
rect 219299 608549 219311 608583
rect 542538 608580 542544 608592
rect 542499 608552 542544 608580
rect 219253 608543 219311 608549
rect 542538 608540 542544 608552
rect 542596 608540 542602 608592
rect 559098 608580 559104 608592
rect 559059 608552 559104 608580
rect 559098 608540 559104 608552
rect 559156 608540 559162 608592
rect 270402 603100 270408 603152
rect 270460 603140 270466 603152
rect 580166 603140 580172 603152
rect 270460 603112 580172 603140
rect 270460 603100 270466 603112
rect 580166 603100 580172 603112
rect 580224 603100 580230 603152
rect 542541 601715 542599 601721
rect 542541 601681 542553 601715
rect 542587 601712 542599 601715
rect 542722 601712 542728 601724
rect 542587 601684 542728 601712
rect 542587 601681 542599 601684
rect 542541 601675 542599 601681
rect 542722 601672 542728 601684
rect 542780 601672 542786 601724
rect 559101 601715 559159 601721
rect 559101 601681 559113 601715
rect 559147 601712 559159 601715
rect 559282 601712 559288 601724
rect 559147 601684 559288 601712
rect 559147 601681 559159 601684
rect 559101 601675 559159 601681
rect 559282 601672 559288 601684
rect 559340 601672 559346 601724
rect 219250 601576 219256 601588
rect 219211 601548 219256 601576
rect 219250 601536 219256 601548
rect 219308 601536 219314 601588
rect 219161 598927 219219 598933
rect 219161 598893 219173 598927
rect 219207 598924 219219 598927
rect 219250 598924 219256 598936
rect 219207 598896 219256 598924
rect 219207 598893 219219 598896
rect 219161 598887 219219 598893
rect 219250 598884 219256 598896
rect 219308 598884 219314 598936
rect 542722 598924 542728 598936
rect 542683 598896 542728 598924
rect 542722 598884 542728 598896
rect 542780 598884 542786 598936
rect 559282 598924 559288 598936
rect 559243 598896 559288 598924
rect 559282 598884 559288 598896
rect 559340 598884 559346 598936
rect 154298 596164 154304 596216
rect 154356 596204 154362 596216
rect 154482 596204 154488 596216
rect 154356 596176 154488 596204
rect 154356 596164 154362 596176
rect 154482 596164 154488 596176
rect 154540 596164 154546 596216
rect 494054 596164 494060 596216
rect 494112 596204 494118 596216
rect 494238 596204 494244 596216
rect 494112 596176 494244 596204
rect 494112 596164 494118 596176
rect 494238 596164 494244 596176
rect 494296 596164 494302 596216
rect 3234 594804 3240 594856
rect 3292 594844 3298 594856
rect 309226 594844 309232 594856
rect 3292 594816 309232 594844
rect 3292 594804 3298 594816
rect 309226 594804 309232 594816
rect 309284 594804 309290 594856
rect 270310 592016 270316 592068
rect 270368 592056 270374 592068
rect 580166 592056 580172 592068
rect 270368 592028 580172 592056
rect 270368 592016 270374 592028
rect 580166 592016 580172 592028
rect 580224 592016 580230 592068
rect 219158 589336 219164 589348
rect 219119 589308 219164 589336
rect 219158 589296 219164 589308
rect 219216 589296 219222 589348
rect 542725 589339 542783 589345
rect 542725 589305 542737 589339
rect 542771 589336 542783 589339
rect 542814 589336 542820 589348
rect 542771 589308 542820 589336
rect 542771 589305 542783 589308
rect 542725 589299 542783 589305
rect 542814 589296 542820 589308
rect 542872 589296 542878 589348
rect 559285 589339 559343 589345
rect 559285 589305 559297 589339
rect 559331 589336 559343 589339
rect 559374 589336 559380 589348
rect 559331 589308 559380 589336
rect 559331 589305 559343 589308
rect 559285 589299 559343 589305
rect 559374 589296 559380 589308
rect 559432 589296 559438 589348
rect 154298 589268 154304 589280
rect 154259 589240 154304 589268
rect 154298 589228 154304 589240
rect 154356 589228 154362 589280
rect 493870 589228 493876 589280
rect 493928 589268 493934 589280
rect 494146 589268 494152 589280
rect 493928 589240 494152 589268
rect 493928 589228 493934 589240
rect 494146 589228 494152 589240
rect 494204 589228 494210 589280
rect 542814 582468 542820 582480
rect 542740 582440 542820 582468
rect 218974 582360 218980 582412
rect 219032 582400 219038 582412
rect 219158 582400 219164 582412
rect 219032 582372 219164 582400
rect 219032 582360 219038 582372
rect 219158 582360 219164 582372
rect 219216 582360 219222 582412
rect 542740 582344 542768 582440
rect 542814 582428 542820 582440
rect 542872 582428 542878 582480
rect 559374 582468 559380 582480
rect 559300 582440 559380 582468
rect 559300 582344 559328 582440
rect 559374 582428 559380 582440
rect 559432 582428 559438 582480
rect 542722 582292 542728 582344
rect 542780 582292 542786 582344
rect 559282 582292 559288 582344
rect 559340 582292 559346 582344
rect 154298 579748 154304 579760
rect 154259 579720 154304 579748
rect 154298 579708 154304 579720
rect 154356 579708 154362 579760
rect 269022 579640 269028 579692
rect 269080 579680 269086 579692
rect 580166 579680 580172 579692
rect 269080 579652 580172 579680
rect 269080 579640 269086 579652
rect 580166 579640 580172 579652
rect 580224 579640 580230 579692
rect 154206 579572 154212 579624
rect 154264 579612 154270 579624
rect 154390 579612 154396 579624
rect 154264 579584 154396 579612
rect 154264 579572 154270 579584
rect 154390 579572 154396 579584
rect 154448 579572 154454 579624
rect 218885 579615 218943 579621
rect 218885 579581 218897 579615
rect 218931 579612 218943 579615
rect 218974 579612 218980 579624
rect 218931 579584 218980 579612
rect 218931 579581 218943 579584
rect 218885 579575 218943 579581
rect 218974 579572 218980 579584
rect 219032 579572 219038 579624
rect 218882 569956 218888 569968
rect 218843 569928 218888 569956
rect 218882 569916 218888 569928
rect 218940 569916 218946 569968
rect 494146 569888 494152 569900
rect 494107 569860 494152 569888
rect 494146 569848 494152 569860
rect 494204 569848 494210 569900
rect 3418 567196 3424 567248
rect 3476 567236 3482 567248
rect 311894 567236 311900 567248
rect 3476 567208 311900 567236
rect 3476 567196 3482 567208
rect 311894 567196 311900 567208
rect 311952 567196 311958 567248
rect 542446 563116 542452 563168
rect 542504 563116 542510 563168
rect 559006 563116 559012 563168
rect 559064 563116 559070 563168
rect 218882 563048 218888 563100
rect 218940 563048 218946 563100
rect 494149 563091 494207 563097
rect 494149 563057 494161 563091
rect 494195 563088 494207 563091
rect 494330 563088 494336 563100
rect 494195 563060 494336 563088
rect 494195 563057 494207 563060
rect 494149 563051 494207 563057
rect 494330 563048 494336 563060
rect 494388 563048 494394 563100
rect 154206 562912 154212 562964
rect 154264 562952 154270 562964
rect 154390 562952 154396 562964
rect 154264 562924 154396 562952
rect 154264 562912 154270 562924
rect 154390 562912 154396 562924
rect 154448 562912 154454 562964
rect 218900 562952 218928 563048
rect 542464 563032 542492 563116
rect 559024 563032 559052 563116
rect 542446 562980 542452 563032
rect 542504 562980 542510 563032
rect 559006 562980 559012 563032
rect 559064 562980 559070 563032
rect 218974 562952 218980 562964
rect 218900 562924 218980 562952
rect 218974 562912 218980 562924
rect 219032 562912 219038 562964
rect 542446 560232 542452 560244
rect 542407 560204 542452 560232
rect 542446 560192 542452 560204
rect 542504 560192 542510 560244
rect 559006 560232 559012 560244
rect 558967 560204 559012 560232
rect 559006 560192 559012 560204
rect 559064 560192 559070 560244
rect 266262 556180 266268 556232
rect 266320 556220 266326 556232
rect 580166 556220 580172 556232
rect 266320 556192 580172 556220
rect 266320 556180 266326 556192
rect 580166 556180 580172 556192
rect 580224 556180 580230 556232
rect 218882 553432 218888 553444
rect 218843 553404 218888 553432
rect 218882 553392 218888 553404
rect 218940 553392 218946 553444
rect 3142 552032 3148 552084
rect 3200 552072 3206 552084
rect 311158 552072 311164 552084
rect 3200 552044 311164 552072
rect 3200 552032 3206 552044
rect 311158 552032 311164 552044
rect 311216 552032 311222 552084
rect 218882 550644 218888 550656
rect 218843 550616 218888 550644
rect 218882 550604 218888 550616
rect 218940 550604 218946 550656
rect 494146 550604 494152 550656
rect 494204 550644 494210 550656
rect 494422 550644 494428 550656
rect 494204 550616 494428 550644
rect 494204 550604 494210 550616
rect 494422 550604 494428 550616
rect 494480 550604 494486 550656
rect 542449 550647 542507 550653
rect 542449 550613 542461 550647
rect 542495 550644 542507 550647
rect 542630 550644 542636 550656
rect 542495 550616 542636 550644
rect 542495 550613 542507 550616
rect 542449 550607 542507 550613
rect 542630 550604 542636 550616
rect 542688 550604 542694 550656
rect 559009 550647 559067 550653
rect 559009 550613 559021 550647
rect 559055 550644 559067 550647
rect 559190 550644 559196 550656
rect 559055 550616 559196 550644
rect 559055 550613 559067 550616
rect 559009 550607 559067 550613
rect 559190 550604 559196 550616
rect 559248 550604 559254 550656
rect 267550 545096 267556 545148
rect 267608 545136 267614 545148
rect 580166 545136 580172 545148
rect 267608 545108 580172 545136
rect 267608 545096 267614 545108
rect 580166 545096 580172 545108
rect 580224 545096 580230 545148
rect 494422 543844 494428 543856
rect 494348 543816 494428 543844
rect 218882 543736 218888 543788
rect 218940 543736 218946 543788
rect 218900 543640 218928 543736
rect 494348 543720 494376 543816
rect 494422 543804 494428 543816
rect 494480 543804 494486 543856
rect 494330 543668 494336 543720
rect 494388 543668 494394 543720
rect 218974 543640 218980 543652
rect 218900 543612 218980 543640
rect 218974 543600 218980 543612
rect 219032 543600 219038 543652
rect 542446 543600 542452 543652
rect 542504 543640 542510 543652
rect 542630 543640 542636 543652
rect 542504 543612 542636 543640
rect 542504 543600 542510 543612
rect 542630 543600 542636 543612
rect 542688 543600 542694 543652
rect 559006 543600 559012 543652
rect 559064 543640 559070 543652
rect 559190 543640 559196 543652
rect 559064 543612 559196 543640
rect 559064 543600 559070 543612
rect 559190 543600 559196 543612
rect 559248 543600 559254 543652
rect 3418 538228 3424 538280
rect 3476 538268 3482 538280
rect 313366 538268 313372 538280
rect 3476 538240 313372 538268
rect 3476 538228 3482 538240
rect 313366 538228 313372 538240
rect 313424 538228 313430 538280
rect 542446 534012 542452 534064
rect 542504 534052 542510 534064
rect 542630 534052 542636 534064
rect 542504 534024 542636 534052
rect 542504 534012 542510 534024
rect 542630 534012 542636 534024
rect 542688 534012 542694 534064
rect 559006 534012 559012 534064
rect 559064 534052 559070 534064
rect 559190 534052 559196 534064
rect 559064 534024 559196 534052
rect 559064 534012 559070 534024
rect 559190 534012 559196 534024
rect 559248 534012 559254 534064
rect 266170 532720 266176 532772
rect 266228 532760 266234 532772
rect 580166 532760 580172 532772
rect 266228 532732 580172 532760
rect 266228 532720 266234 532732
rect 580166 532720 580172 532732
rect 580224 532720 580230 532772
rect 494146 531292 494152 531344
rect 494204 531332 494210 531344
rect 494422 531332 494428 531344
rect 494204 531304 494428 531332
rect 494204 531292 494210 531304
rect 494422 531292 494428 531304
rect 494480 531292 494486 531344
rect 154390 531264 154396 531276
rect 154351 531236 154396 531264
rect 154390 531224 154396 531236
rect 154448 531224 154454 531276
rect 494422 524532 494428 524544
rect 494348 524504 494428 524532
rect 494348 524408 494376 524504
rect 494422 524492 494428 524504
rect 494480 524492 494486 524544
rect 542630 524424 542636 524476
rect 542688 524424 542694 524476
rect 559190 524424 559196 524476
rect 559248 524424 559254 524476
rect 494330 524356 494336 524408
rect 494388 524356 494394 524408
rect 542648 524396 542676 524424
rect 542722 524396 542728 524408
rect 542648 524368 542728 524396
rect 542722 524356 542728 524368
rect 542780 524356 542786 524408
rect 559208 524396 559236 524424
rect 559282 524396 559288 524408
rect 559208 524368 559288 524396
rect 559282 524356 559288 524368
rect 559340 524356 559346 524408
rect 218974 524288 218980 524340
rect 219032 524328 219038 524340
rect 219158 524328 219164 524340
rect 219032 524300 219164 524328
rect 219032 524288 219038 524300
rect 219158 524288 219164 524300
rect 219216 524288 219222 524340
rect 154393 521679 154451 521685
rect 154393 521645 154405 521679
rect 154439 521676 154451 521679
rect 154482 521676 154488 521688
rect 154439 521648 154488 521676
rect 154439 521645 154451 521648
rect 154393 521639 154451 521645
rect 154482 521636 154488 521648
rect 154540 521636 154546 521688
rect 218790 514632 218796 514684
rect 218848 514672 218854 514684
rect 219066 514672 219072 514684
rect 218848 514644 219072 514672
rect 218848 514632 218854 514644
rect 219066 514632 219072 514644
rect 219124 514632 219130 514684
rect 494146 511980 494152 512032
rect 494204 512020 494210 512032
rect 494422 512020 494428 512032
rect 494204 511992 494428 512020
rect 494204 511980 494210 511992
rect 494422 511980 494428 511992
rect 494480 511980 494486 512032
rect 542538 511980 542544 512032
rect 542596 512020 542602 512032
rect 542814 512020 542820 512032
rect 542596 511992 542820 512020
rect 542596 511980 542602 511992
rect 542814 511980 542820 511992
rect 542872 511980 542878 512032
rect 559098 511980 559104 512032
rect 559156 512020 559162 512032
rect 559374 512020 559380 512032
rect 559156 511992 559380 512020
rect 559156 511980 559162 511992
rect 559374 511980 559380 511992
rect 559432 511980 559438 512032
rect 154390 511952 154396 511964
rect 154351 511924 154396 511952
rect 154390 511912 154396 511924
rect 154448 511912 154454 511964
rect 219066 510592 219072 510604
rect 219027 510564 219072 510592
rect 219066 510552 219072 510564
rect 219124 510552 219130 510604
rect 3418 509328 3424 509380
rect 3476 509368 3482 509380
rect 314654 509368 314660 509380
rect 3476 509340 314660 509368
rect 3476 509328 3482 509340
rect 314654 509328 314660 509340
rect 314712 509328 314718 509380
rect 263502 509260 263508 509312
rect 263560 509300 263566 509312
rect 580166 509300 580172 509312
rect 263560 509272 580172 509300
rect 263560 509260 263566 509272
rect 580166 509260 580172 509272
rect 580224 509260 580230 509312
rect 219066 505084 219072 505096
rect 219027 505056 219072 505084
rect 219066 505044 219072 505056
rect 219124 505044 219130 505096
rect 154393 502367 154451 502373
rect 154393 502333 154405 502367
rect 154439 502364 154451 502367
rect 154482 502364 154488 502376
rect 154439 502336 154488 502364
rect 154439 502333 154451 502336
rect 154393 502327 154451 502333
rect 154482 502324 154488 502336
rect 154540 502324 154546 502376
rect 494238 502324 494244 502376
rect 494296 502364 494302 502376
rect 494422 502364 494428 502376
rect 494296 502336 494428 502364
rect 494296 502324 494302 502336
rect 494422 502324 494428 502336
rect 494480 502324 494486 502376
rect 542630 502324 542636 502376
rect 542688 502364 542694 502376
rect 542814 502364 542820 502376
rect 542688 502336 542820 502364
rect 542688 502324 542694 502336
rect 542814 502324 542820 502336
rect 542872 502324 542878 502376
rect 559190 502324 559196 502376
rect 559248 502364 559254 502376
rect 559374 502364 559380 502376
rect 559248 502336 559380 502364
rect 559248 502324 559254 502336
rect 559374 502324 559380 502336
rect 559432 502324 559438 502376
rect 264882 498176 264888 498228
rect 264940 498216 264946 498228
rect 580166 498216 580172 498228
rect 264940 498188 580172 498216
rect 264940 498176 264946 498188
rect 580166 498176 580172 498188
rect 580224 498176 580230 498228
rect 3418 495456 3424 495508
rect 3476 495496 3482 495508
rect 313918 495496 313924 495508
rect 3476 495468 313924 495496
rect 3476 495456 3482 495468
rect 313918 495456 313924 495468
rect 313976 495456 313982 495508
rect 219066 492668 219072 492720
rect 219124 492708 219130 492720
rect 219158 492708 219164 492720
rect 219124 492680 219164 492708
rect 219124 492668 219130 492680
rect 219158 492668 219164 492680
rect 219216 492668 219222 492720
rect 542538 492640 542544 492652
rect 542499 492612 542544 492640
rect 542538 492600 542544 492612
rect 542596 492600 542602 492652
rect 559098 492640 559104 492652
rect 559059 492612 559104 492640
rect 559098 492600 559104 492612
rect 559156 492600 559162 492652
rect 154298 485800 154304 485852
rect 154356 485800 154362 485852
rect 219158 485800 219164 485852
rect 219216 485800 219222 485852
rect 262122 485800 262128 485852
rect 262180 485840 262186 485852
rect 580166 485840 580172 485852
rect 262180 485812 580172 485840
rect 262180 485800 262186 485812
rect 580166 485800 580172 485812
rect 580224 485800 580230 485852
rect 154316 485704 154344 485800
rect 154390 485704 154396 485716
rect 154316 485676 154396 485704
rect 154390 485664 154396 485676
rect 154448 485664 154454 485716
rect 219176 485704 219204 485800
rect 542538 485772 542544 485784
rect 542499 485744 542544 485772
rect 542538 485732 542544 485744
rect 542596 485732 542602 485784
rect 559098 485772 559104 485784
rect 559059 485744 559104 485772
rect 559098 485732 559104 485744
rect 559156 485732 559162 485784
rect 219250 485704 219256 485716
rect 219176 485676 219256 485704
rect 219250 485664 219256 485676
rect 219308 485664 219314 485716
rect 154390 482984 154396 482996
rect 154351 482956 154396 482984
rect 154390 482944 154396 482956
rect 154448 482944 154454 482996
rect 3142 480224 3148 480276
rect 3200 480264 3206 480276
rect 316034 480264 316040 480276
rect 3200 480236 316040 480264
rect 3200 480224 3206 480236
rect 316034 480224 316040 480236
rect 316092 480224 316098 480276
rect 494054 480224 494060 480276
rect 494112 480264 494118 480276
rect 494238 480264 494244 480276
rect 494112 480236 494244 480264
rect 494112 480224 494118 480236
rect 494238 480224 494244 480236
rect 494296 480224 494302 480276
rect 219066 476076 219072 476128
rect 219124 476116 219130 476128
rect 219250 476116 219256 476128
rect 219124 476088 219256 476116
rect 219124 476076 219130 476088
rect 219250 476076 219256 476088
rect 219308 476076 219314 476128
rect 542446 476076 542452 476128
rect 542504 476116 542510 476128
rect 542630 476116 542636 476128
rect 542504 476088 542636 476116
rect 542504 476076 542510 476088
rect 542630 476076 542636 476088
rect 542688 476076 542694 476128
rect 559006 476076 559012 476128
rect 559064 476116 559070 476128
rect 559190 476116 559196 476128
rect 559064 476088 559196 476116
rect 559064 476076 559070 476088
rect 559190 476076 559196 476088
rect 559248 476076 559254 476128
rect 154390 476048 154396 476060
rect 154351 476020 154396 476048
rect 154390 476008 154396 476020
rect 154448 476008 154454 476060
rect 542541 466531 542599 466537
rect 542541 466497 542553 466531
rect 542587 466528 542599 466531
rect 542630 466528 542636 466540
rect 542587 466500 542636 466528
rect 542587 466497 542599 466500
rect 542541 466491 542599 466497
rect 542630 466488 542636 466500
rect 542688 466488 542694 466540
rect 559101 466531 559159 466537
rect 559101 466497 559113 466531
rect 559147 466528 559159 466531
rect 559190 466528 559196 466540
rect 559147 466500 559196 466528
rect 559147 466497 559159 466500
rect 559101 466491 559159 466497
rect 559190 466488 559196 466500
rect 559248 466488 559254 466540
rect 542538 463740 542544 463752
rect 542499 463712 542544 463740
rect 542538 463700 542544 463712
rect 542596 463700 542602 463752
rect 559098 463740 559104 463752
rect 559059 463712 559104 463740
rect 559098 463700 559104 463712
rect 559156 463700 559162 463752
rect 286965 463675 287023 463681
rect 286965 463641 286977 463675
rect 287011 463672 287023 463675
rect 291378 463672 291384 463684
rect 287011 463644 291384 463672
rect 287011 463641 287023 463644
rect 286965 463635 287023 463641
rect 291378 463632 291384 463644
rect 291436 463632 291442 463684
rect 291838 463632 291844 463684
rect 291896 463672 291902 463684
rect 294506 463672 294512 463684
rect 291896 463644 294512 463672
rect 291896 463632 291902 463644
rect 294506 463632 294512 463644
rect 294564 463632 294570 463684
rect 297358 463632 297364 463684
rect 297416 463672 297422 463684
rect 300854 463672 300860 463684
rect 297416 463644 300860 463672
rect 297416 463632 297422 463644
rect 300854 463632 300860 463644
rect 300912 463632 300918 463684
rect 301498 463632 301504 463684
rect 301556 463672 301562 463684
rect 303982 463672 303988 463684
rect 301556 463644 303988 463672
rect 301556 463632 301562 463644
rect 303982 463632 303988 463644
rect 304040 463632 304046 463684
rect 308398 463632 308404 463684
rect 308456 463672 308462 463684
rect 311342 463672 311348 463684
rect 308456 463644 311348 463672
rect 308456 463632 308462 463644
rect 311342 463632 311348 463644
rect 311400 463632 311406 463684
rect 282917 463607 282975 463613
rect 282917 463573 282929 463607
rect 282963 463604 282975 463607
rect 287793 463607 287851 463613
rect 287793 463604 287805 463607
rect 282963 463576 287805 463604
rect 282963 463573 282975 463576
rect 282917 463567 282975 463573
rect 287793 463573 287805 463576
rect 287839 463573 287851 463607
rect 287793 463567 287851 463573
rect 290458 463564 290464 463616
rect 290516 463604 290522 463616
rect 293494 463604 293500 463616
rect 290516 463576 293500 463604
rect 290516 463564 290522 463576
rect 293494 463564 293500 463576
rect 293552 463564 293558 463616
rect 293589 463607 293647 463613
rect 293589 463573 293601 463607
rect 293635 463604 293647 463607
rect 298738 463604 298744 463616
rect 293635 463576 298744 463604
rect 293635 463573 293647 463576
rect 293589 463567 293647 463573
rect 298738 463564 298744 463576
rect 298796 463564 298802 463616
rect 300118 463564 300124 463616
rect 300176 463604 300182 463616
rect 302970 463604 302976 463616
rect 300176 463576 302976 463604
rect 300176 463564 300182 463576
rect 302970 463564 302976 463576
rect 303028 463564 303034 463616
rect 311158 463564 311164 463616
rect 311216 463604 311222 463616
rect 314562 463604 314568 463616
rect 311216 463576 314568 463604
rect 311216 463564 311222 463576
rect 314562 463564 314568 463576
rect 314620 463564 314626 463616
rect 259457 463539 259515 463545
rect 259457 463505 259469 463539
rect 259503 463536 259515 463539
rect 269025 463539 269083 463545
rect 269025 463536 269037 463539
rect 259503 463508 269037 463536
rect 259503 463505 259515 463508
rect 259457 463499 259515 463505
rect 269025 463505 269037 463508
rect 269071 463505 269083 463539
rect 269025 463499 269083 463505
rect 269117 463539 269175 463545
rect 269117 463505 269129 463539
rect 269163 463536 269175 463539
rect 278685 463539 278743 463545
rect 278685 463536 278697 463539
rect 269163 463508 278697 463536
rect 269163 463505 269175 463508
rect 269117 463499 269175 463505
rect 278685 463505 278697 463508
rect 278731 463505 278743 463539
rect 278685 463499 278743 463505
rect 280890 463496 280896 463548
rect 280948 463536 280954 463548
rect 287057 463539 287115 463545
rect 287057 463536 287069 463539
rect 280948 463508 287069 463536
rect 280948 463496 280954 463508
rect 287057 463505 287069 463508
rect 287103 463505 287115 463539
rect 287057 463499 287115 463505
rect 287701 463539 287759 463545
rect 287701 463505 287713 463539
rect 287747 463536 287759 463539
rect 296625 463539 296683 463545
rect 296625 463536 296637 463539
rect 287747 463508 296637 463536
rect 287747 463505 287759 463508
rect 287701 463499 287759 463505
rect 296625 463505 296637 463508
rect 296671 463505 296683 463539
rect 296625 463499 296683 463505
rect 267642 463428 267648 463480
rect 267700 463468 267706 463480
rect 286965 463471 287023 463477
rect 286965 463468 286977 463471
rect 267700 463440 286977 463468
rect 267700 463428 267706 463440
rect 286965 463437 286977 463440
rect 287011 463437 287023 463471
rect 286965 463431 287023 463437
rect 287241 463471 287299 463477
rect 287241 463437 287253 463471
rect 287287 463468 287299 463471
rect 291197 463471 291255 463477
rect 291197 463468 291209 463471
rect 287287 463440 291209 463468
rect 287287 463437 287299 463440
rect 287241 463431 287299 463437
rect 291197 463437 291209 463440
rect 291243 463437 291255 463471
rect 291197 463431 291255 463437
rect 291289 463471 291347 463477
rect 291289 463437 291301 463471
rect 291335 463468 291347 463471
rect 295610 463468 295616 463480
rect 291335 463440 295616 463468
rect 291335 463437 291347 463440
rect 291289 463431 291347 463437
rect 295610 463428 295616 463440
rect 295668 463428 295674 463480
rect 295978 463428 295984 463480
rect 296036 463468 296042 463480
rect 299750 463468 299756 463480
rect 296036 463440 299756 463468
rect 296036 463428 296042 463440
rect 299750 463428 299756 463440
rect 299808 463428 299814 463480
rect 96617 463403 96675 463409
rect 96617 463369 96629 463403
rect 96663 463400 96675 463403
rect 106185 463403 106243 463409
rect 106185 463400 106197 463403
rect 96663 463372 106197 463400
rect 96663 463369 96675 463372
rect 96617 463363 96675 463369
rect 106185 463369 106197 463372
rect 106231 463369 106243 463403
rect 106185 463363 106243 463369
rect 157337 463403 157395 463409
rect 157337 463369 157349 463403
rect 157383 463400 157395 463403
rect 160925 463403 160983 463409
rect 160925 463400 160937 463403
rect 157383 463372 160937 463400
rect 157383 463369 157395 463372
rect 157337 463363 157395 463369
rect 160925 463369 160937 463372
rect 160971 463369 160983 463403
rect 160925 463363 160983 463369
rect 183557 463403 183615 463409
rect 183557 463369 183569 463403
rect 183603 463400 183615 463403
rect 193125 463403 193183 463409
rect 193125 463400 193137 463403
rect 183603 463372 193137 463400
rect 183603 463369 183615 463372
rect 183557 463363 183615 463369
rect 193125 463369 193137 463372
rect 193171 463369 193183 463403
rect 193125 463363 193183 463369
rect 200117 463403 200175 463409
rect 200117 463369 200129 463403
rect 200163 463400 200175 463403
rect 205637 463403 205695 463409
rect 205637 463400 205649 463403
rect 200163 463372 205649 463400
rect 200163 463369 200175 463372
rect 200117 463363 200175 463369
rect 205637 463369 205649 463372
rect 205683 463369 205695 463403
rect 205637 463363 205695 463369
rect 219066 463360 219072 463412
rect 219124 463400 219130 463412
rect 282917 463403 282975 463409
rect 282917 463400 282929 463403
rect 219124 463372 282929 463400
rect 219124 463360 219130 463372
rect 282917 463369 282929 463372
rect 282963 463369 282975 463403
rect 282917 463363 282975 463369
rect 283009 463403 283067 463409
rect 283009 463369 283021 463403
rect 283055 463400 283067 463403
rect 287701 463403 287759 463409
rect 287701 463400 287713 463403
rect 283055 463372 287713 463400
rect 283055 463369 283067 463372
rect 283009 463363 283067 463369
rect 287701 463369 287713 463372
rect 287747 463369 287759 463403
rect 287701 463363 287759 463369
rect 293218 463360 293224 463412
rect 293276 463400 293282 463412
rect 296622 463400 296628 463412
rect 293276 463372 296628 463400
rect 293276 463360 293282 463372
rect 296622 463360 296628 463372
rect 296680 463360 296686 463412
rect 125597 463335 125655 463341
rect 125597 463301 125609 463335
rect 125643 463332 125655 463335
rect 129734 463332 129740 463344
rect 125643 463304 129740 463332
rect 125643 463301 125655 463304
rect 125597 463295 125655 463301
rect 129734 463292 129740 463304
rect 129792 463292 129798 463344
rect 154298 463292 154304 463344
rect 154356 463332 154362 463344
rect 293589 463335 293647 463341
rect 293589 463332 293601 463335
rect 154356 463304 293601 463332
rect 154356 463292 154362 463304
rect 293589 463301 293601 463304
rect 293635 463301 293647 463335
rect 293589 463295 293647 463301
rect 294598 463292 294604 463344
rect 294656 463332 294662 463344
rect 297726 463332 297732 463344
rect 294656 463304 297732 463332
rect 294656 463292 294662 463304
rect 297726 463292 297732 463304
rect 297784 463292 297790 463344
rect 89717 463267 89775 463273
rect 89717 463233 89729 463267
rect 89763 463264 89775 463267
rect 96617 463267 96675 463273
rect 96617 463264 96629 463267
rect 89763 463236 96629 463264
rect 89763 463233 89775 463236
rect 89717 463227 89775 463233
rect 96617 463233 96629 463236
rect 96663 463233 96675 463267
rect 96617 463227 96675 463233
rect 129826 463224 129832 463276
rect 129884 463264 129890 463276
rect 160925 463267 160983 463273
rect 129884 463236 138244 463264
rect 129884 463224 129890 463236
rect 106185 463199 106243 463205
rect 106185 463165 106197 463199
rect 106231 463196 106243 463199
rect 125597 463199 125655 463205
rect 125597 463196 125609 463199
rect 106231 463168 108988 463196
rect 106231 463165 106243 463168
rect 106185 463159 106243 463165
rect 89622 463088 89628 463140
rect 89680 463128 89686 463140
rect 89717 463131 89775 463137
rect 89717 463128 89729 463131
rect 89680 463100 89729 463128
rect 89680 463088 89686 463100
rect 89717 463097 89729 463100
rect 89763 463097 89775 463131
rect 108960 463128 108988 463168
rect 120644 463168 125609 463196
rect 118605 463131 118663 463137
rect 118605 463128 118617 463131
rect 108960 463100 118617 463128
rect 89717 463091 89775 463097
rect 118605 463097 118617 463100
rect 118651 463097 118663 463131
rect 118605 463091 118663 463097
rect 118697 463131 118755 463137
rect 118697 463097 118709 463131
rect 118743 463128 118755 463131
rect 120644 463128 120672 463168
rect 125597 463165 125609 463168
rect 125643 463165 125655 463199
rect 138216 463196 138244 463236
rect 160925 463233 160937 463267
rect 160971 463264 160983 463267
rect 173897 463267 173955 463273
rect 173897 463264 173909 463267
rect 160971 463236 173909 463264
rect 160971 463233 160983 463236
rect 160925 463227 160983 463233
rect 173897 463233 173909 463236
rect 173943 463233 173955 463267
rect 173897 463227 173955 463233
rect 195885 463267 195943 463273
rect 195885 463233 195897 463267
rect 195931 463264 195943 463267
rect 269117 463267 269175 463273
rect 195931 463236 196480 463264
rect 195931 463233 195943 463236
rect 195885 463227 195943 463233
rect 147674 463196 147680 463208
rect 138216 463168 147680 463196
rect 125597 463159 125655 463165
rect 147674 463156 147680 463168
rect 147732 463156 147738 463208
rect 183465 463199 183523 463205
rect 183465 463165 183477 463199
rect 183511 463165 183523 463199
rect 183465 463159 183523 463165
rect 183557 463199 183615 463205
rect 183557 463165 183569 463199
rect 183603 463165 183615 463199
rect 183557 463159 183615 463165
rect 193125 463199 193183 463205
rect 193125 463165 193137 463199
rect 193171 463196 193183 463199
rect 195793 463199 195851 463205
rect 195793 463196 195805 463199
rect 193171 463168 195805 463196
rect 193171 463165 193183 463168
rect 193125 463159 193183 463165
rect 195793 463165 195805 463168
rect 195839 463165 195851 463199
rect 196452 463196 196480 463236
rect 209884 463236 215432 463264
rect 200117 463199 200175 463205
rect 200117 463196 200129 463199
rect 196452 463168 200129 463196
rect 195793 463159 195851 463165
rect 200117 463165 200129 463168
rect 200163 463165 200175 463199
rect 200117 463159 200175 463165
rect 205637 463199 205695 463205
rect 205637 463165 205649 463199
rect 205683 463196 205695 463199
rect 209884 463196 209912 463236
rect 205683 463168 209912 463196
rect 215404 463196 215432 463236
rect 269117 463233 269129 463267
rect 269163 463233 269175 463267
rect 269117 463227 269175 463233
rect 278685 463267 278743 463273
rect 278685 463233 278697 463267
rect 278731 463264 278743 463267
rect 283009 463267 283067 463273
rect 283009 463264 283021 463267
rect 278731 463236 283021 463264
rect 278731 463233 278743 463236
rect 278685 463227 278743 463233
rect 283009 463233 283021 463236
rect 283055 463233 283067 463267
rect 283009 463227 283067 463233
rect 287793 463267 287851 463273
rect 287793 463233 287805 463267
rect 287839 463264 287851 463267
rect 291289 463267 291347 463273
rect 291289 463264 291301 463267
rect 287839 463236 291301 463264
rect 287839 463233 287851 463236
rect 287793 463227 287851 463233
rect 291289 463233 291301 463236
rect 291335 463233 291347 463267
rect 291289 463227 291347 463233
rect 296625 463267 296683 463273
rect 296625 463233 296637 463267
rect 296671 463264 296683 463267
rect 301866 463264 301872 463276
rect 296671 463236 301872 463264
rect 296671 463233 296683 463236
rect 296625 463227 296683 463233
rect 222197 463199 222255 463205
rect 222197 463196 222209 463199
rect 215404 463168 222209 463196
rect 205683 463165 205695 463168
rect 205637 463159 205695 463165
rect 222197 463165 222209 463168
rect 222243 463165 222255 463199
rect 222197 463159 222255 463165
rect 222289 463199 222347 463205
rect 222289 463165 222301 463199
rect 222335 463196 222347 463199
rect 234525 463199 234583 463205
rect 234525 463196 234537 463199
rect 222335 463168 234537 463196
rect 222335 463165 222347 463168
rect 222289 463159 222347 463165
rect 234525 463165 234537 463168
rect 234571 463165 234583 463199
rect 234525 463159 234583 463165
rect 234617 463199 234675 463205
rect 234617 463165 234629 463199
rect 234663 463196 234675 463199
rect 244185 463199 244243 463205
rect 244185 463196 244197 463199
rect 234663 463168 244197 463196
rect 234663 463165 234675 463168
rect 234617 463159 234675 463165
rect 244185 463165 244197 463168
rect 244231 463165 244243 463199
rect 244185 463159 244243 463165
rect 244277 463199 244335 463205
rect 244277 463165 244289 463199
rect 244323 463196 244335 463199
rect 253845 463199 253903 463205
rect 253845 463196 253857 463199
rect 244323 463168 253857 463196
rect 244323 463165 244335 463168
rect 244277 463159 244335 463165
rect 253845 463165 253857 463168
rect 253891 463165 253903 463199
rect 253845 463159 253903 463165
rect 253937 463199 253995 463205
rect 253937 463165 253949 463199
rect 253983 463196 253995 463199
rect 259457 463199 259515 463205
rect 259457 463196 259469 463199
rect 253983 463168 259469 463196
rect 253983 463165 253995 463168
rect 253937 463159 253995 463165
rect 259457 463165 259469 463168
rect 259503 463165 259515 463199
rect 259457 463159 259515 463165
rect 269025 463199 269083 463205
rect 269025 463165 269037 463199
rect 269071 463196 269083 463199
rect 269132 463196 269160 463227
rect 301866 463224 301872 463236
rect 301924 463224 301930 463276
rect 269071 463168 269160 463196
rect 269071 463165 269083 463168
rect 269025 463159 269083 463165
rect 118743 463100 120672 463128
rect 118743 463097 118755 463100
rect 118697 463091 118755 463097
rect 147766 463088 147772 463140
rect 147824 463128 147830 463140
rect 157337 463131 157395 463137
rect 157337 463128 157349 463131
rect 147824 463100 157349 463128
rect 147824 463088 147830 463100
rect 157337 463097 157349 463100
rect 157383 463097 157395 463131
rect 183480 463128 183508 463159
rect 183572 463128 183600 463159
rect 279786 463156 279792 463208
rect 279844 463196 279850 463208
rect 279844 463168 280292 463196
rect 279844 463156 279850 463168
rect 183480 463100 183600 463128
rect 157337 463091 157395 463097
rect 277670 463088 277676 463140
rect 277728 463128 277734 463140
rect 280264 463128 280292 463168
rect 281902 463156 281908 463208
rect 281960 463196 281966 463208
rect 282822 463196 282828 463208
rect 281960 463168 282828 463196
rect 281960 463156 281966 463168
rect 282822 463156 282828 463168
rect 282880 463156 282886 463208
rect 282914 463156 282920 463208
rect 282972 463196 282978 463208
rect 284110 463196 284116 463208
rect 282972 463168 284116 463196
rect 282972 463156 282978 463168
rect 284110 463156 284116 463168
rect 284168 463156 284174 463208
rect 286134 463156 286140 463208
rect 286192 463196 286198 463208
rect 286962 463196 286968 463208
rect 286192 463168 286968 463196
rect 286192 463156 286198 463168
rect 286962 463156 286968 463168
rect 287020 463156 287026 463208
rect 287146 463156 287152 463208
rect 287204 463196 287210 463208
rect 288342 463196 288348 463208
rect 287204 463168 288348 463196
rect 287204 463156 287210 463168
rect 288342 463156 288348 463168
rect 288400 463156 288406 463208
rect 290366 463156 290372 463208
rect 290424 463196 290430 463208
rect 291102 463196 291108 463208
rect 290424 463168 291108 463196
rect 290424 463156 290430 463168
rect 291102 463156 291108 463168
rect 291160 463156 291166 463208
rect 291197 463199 291255 463205
rect 291197 463165 291209 463199
rect 291243 463196 291255 463199
rect 494238 463196 494244 463208
rect 291243 463168 494244 463196
rect 291243 463165 291255 463168
rect 291197 463159 291255 463165
rect 494238 463156 494244 463168
rect 494296 463156 494302 463208
rect 542538 463128 542544 463140
rect 277728 463100 280200 463128
rect 280264 463100 542544 463128
rect 277728 463088 277734 463100
rect 24762 463020 24768 463072
rect 24820 463060 24826 463072
rect 279973 463063 280031 463069
rect 279973 463060 279985 463063
rect 24820 463032 279985 463060
rect 24820 463020 24826 463032
rect 279973 463029 279985 463032
rect 280019 463029 280031 463063
rect 279973 463023 280031 463029
rect 173897 462995 173955 463001
rect 173897 462961 173909 462995
rect 173943 462992 173955 462995
rect 183465 462995 183523 463001
rect 183465 462992 183477 462995
rect 173943 462964 183477 462992
rect 173943 462961 173955 462964
rect 173897 462955 173955 462961
rect 183465 462961 183477 462964
rect 183511 462961 183523 462995
rect 183465 462955 183523 462961
rect 264054 462952 264060 463004
rect 264112 462992 264118 463004
rect 264882 462992 264888 463004
rect 264112 462964 264888 462992
rect 264112 462952 264118 462964
rect 264882 462952 264888 462964
rect 264940 462952 264946 463004
rect 265066 462952 265072 463004
rect 265124 462992 265130 463004
rect 266170 462992 266176 463004
rect 265124 462964 266176 462992
rect 265124 462952 265130 462964
rect 266170 462952 266176 462964
rect 266228 462952 266234 463004
rect 268194 462952 268200 463004
rect 268252 462992 268258 463004
rect 269022 462992 269028 463004
rect 268252 462964 269028 462992
rect 268252 462952 268258 462964
rect 269022 462952 269028 462964
rect 269080 462952 269086 463004
rect 269298 462952 269304 463004
rect 269356 462992 269362 463004
rect 270402 462992 270408 463004
rect 269356 462964 270408 462992
rect 269356 462952 269362 462964
rect 270402 462952 270408 462964
rect 270460 462952 270466 463004
rect 272426 462952 272432 463004
rect 272484 462992 272490 463004
rect 273162 462992 273168 463004
rect 272484 462964 273168 462992
rect 272484 462952 272490 462964
rect 273162 462952 273168 462964
rect 273220 462952 273226 463004
rect 273438 462952 273444 463004
rect 273496 462992 273502 463004
rect 274450 462992 274456 463004
rect 273496 462964 274456 462992
rect 273496 462952 273502 462964
rect 274450 462952 274456 462964
rect 274508 462952 274514 463004
rect 278774 462952 278780 463004
rect 278832 462992 278838 463004
rect 280062 462992 280068 463004
rect 278832 462964 280068 462992
rect 278832 462952 278838 462964
rect 280062 462952 280068 462964
rect 280120 462952 280126 463004
rect 280172 462992 280200 463100
rect 542538 463088 542544 463100
rect 542596 463088 542602 463140
rect 280249 463063 280307 463069
rect 280249 463029 280261 463063
rect 280295 463060 280307 463063
rect 304994 463060 305000 463072
rect 280295 463032 305000 463060
rect 280295 463029 280307 463032
rect 280249 463023 280307 463029
rect 304994 463020 305000 463032
rect 305052 463020 305058 463072
rect 305638 463020 305644 463072
rect 305696 463060 305702 463072
rect 308214 463060 308220 463072
rect 305696 463032 308220 463060
rect 305696 463020 305702 463032
rect 308214 463020 308220 463032
rect 308272 463020 308278 463072
rect 313918 463020 313924 463072
rect 313976 463060 313982 463072
rect 317690 463060 317696 463072
rect 313976 463032 317696 463060
rect 313976 463020 313982 463032
rect 317690 463020 317696 463032
rect 317748 463020 317754 463072
rect 559098 462992 559104 463004
rect 280172 462964 559104 462992
rect 559098 462952 559104 462964
rect 559156 462952 559162 463004
rect 31018 462884 31024 462936
rect 31076 462924 31082 462936
rect 342898 462924 342904 462936
rect 31076 462896 342904 462924
rect 31076 462884 31082 462896
rect 342898 462884 342904 462896
rect 342956 462884 342962 462936
rect 4614 462816 4620 462868
rect 4672 462856 4678 462868
rect 320818 462856 320824 462868
rect 4672 462828 320824 462856
rect 4672 462816 4678 462828
rect 320818 462816 320824 462828
rect 320876 462816 320882 462868
rect 2958 462748 2964 462800
rect 3016 462788 3022 462800
rect 319806 462788 319812 462800
rect 3016 462760 319812 462788
rect 3016 462748 3022 462760
rect 319806 462748 319812 462760
rect 319864 462748 319870 462800
rect 3234 462680 3240 462732
rect 3292 462720 3298 462732
rect 322934 462720 322940 462732
rect 3292 462692 322940 462720
rect 3292 462680 3298 462692
rect 322934 462680 322940 462692
rect 322992 462680 322998 462732
rect 3142 462612 3148 462664
rect 3200 462652 3206 462664
rect 324038 462652 324044 462664
rect 3200 462624 324044 462652
rect 3200 462612 3206 462624
rect 324038 462612 324044 462624
rect 324096 462612 324102 462664
rect 259822 462544 259828 462596
rect 259880 462584 259886 462596
rect 580074 462584 580080 462596
rect 259880 462556 580080 462584
rect 259880 462544 259886 462556
rect 580074 462544 580080 462556
rect 580132 462544 580138 462596
rect 238754 462476 238760 462528
rect 238812 462516 238818 462528
rect 577498 462516 577504 462528
rect 238812 462488 577504 462516
rect 238812 462476 238818 462488
rect 577498 462476 577504 462488
rect 577556 462476 577562 462528
rect 236638 462408 236644 462460
rect 236696 462448 236702 462460
rect 580350 462448 580356 462460
rect 236696 462420 580356 462448
rect 236696 462408 236702 462420
rect 580350 462408 580356 462420
rect 580408 462408 580414 462460
rect 3418 462340 3424 462392
rect 3476 462380 3482 462392
rect 348234 462380 348240 462392
rect 3476 462352 348240 462380
rect 3476 462340 3482 462352
rect 348234 462340 348240 462352
rect 348292 462340 348298 462392
rect 260834 460232 260840 460284
rect 260892 460272 260898 460284
rect 580166 460272 580172 460284
rect 260892 460244 580172 460272
rect 260892 460232 260898 460244
rect 580166 460232 580172 460244
rect 580224 460232 580230 460284
rect 4706 460164 4712 460216
rect 4764 460204 4770 460216
rect 327166 460204 327172 460216
rect 4764 460176 327172 460204
rect 4764 460164 4770 460176
rect 327166 460164 327172 460176
rect 327224 460164 327230 460216
rect 5442 460096 5448 460148
rect 5500 460136 5506 460148
rect 330294 460136 330300 460148
rect 5500 460108 330300 460136
rect 5500 460096 5506 460108
rect 330294 460096 330300 460108
rect 330352 460096 330358 460148
rect 5258 460028 5264 460080
rect 5316 460068 5322 460080
rect 333054 460068 333060 460080
rect 5316 460040 333060 460068
rect 5316 460028 5322 460040
rect 333054 460028 333060 460040
rect 333112 460028 333118 460080
rect 250714 459960 250720 460012
rect 250772 460000 250778 460012
rect 579982 460000 579988 460012
rect 250772 459972 579988 460000
rect 250772 459960 250778 459972
rect 579982 459960 579988 459972
rect 580040 459960 580046 460012
rect 5074 459892 5080 459944
rect 5132 459932 5138 459944
rect 336366 459932 336372 459944
rect 5132 459904 336372 459932
rect 5132 459892 5138 459904
rect 336366 459892 336372 459904
rect 336424 459892 336430 459944
rect 247586 459824 247592 459876
rect 247644 459864 247650 459876
rect 579706 459864 579712 459876
rect 247644 459836 579712 459864
rect 247644 459824 247650 459836
rect 579706 459824 579712 459836
rect 579764 459824 579770 459876
rect 4890 459756 4896 459808
rect 4948 459796 4954 459808
rect 339494 459796 339500 459808
rect 4948 459768 339500 459796
rect 4948 459756 4954 459768
rect 339494 459756 339500 459768
rect 339552 459756 339558 459808
rect 244090 459688 244096 459740
rect 244148 459728 244154 459740
rect 580810 459728 580816 459740
rect 244148 459700 580816 459728
rect 244148 459688 244154 459700
rect 580810 459688 580816 459700
rect 580868 459688 580874 459740
rect 241146 459620 241152 459672
rect 241204 459660 241210 459672
rect 580626 459660 580632 459672
rect 241204 459632 580632 459660
rect 241204 459620 241210 459632
rect 580626 459620 580632 459632
rect 580684 459620 580690 459672
rect 235902 459552 235908 459604
rect 235960 459592 235966 459604
rect 580258 459592 580264 459604
rect 235960 459564 580264 459592
rect 235960 459552 235966 459564
rect 580258 459552 580264 459564
rect 580316 459552 580322 459604
rect 247405 459527 247463 459533
rect 247405 459493 247417 459527
rect 247451 459524 247463 459527
rect 258721 459527 258779 459533
rect 258721 459524 258733 459527
rect 247451 459496 258733 459524
rect 247451 459493 247463 459496
rect 247405 459487 247463 459493
rect 258721 459493 258733 459496
rect 258767 459493 258779 459527
rect 258721 459487 258779 459493
rect 268381 459527 268439 459533
rect 268381 459493 268393 459527
rect 268427 459524 268439 459527
rect 278041 459527 278099 459533
rect 278041 459524 278053 459527
rect 268427 459496 278053 459524
rect 268427 459493 268439 459496
rect 268381 459487 268439 459493
rect 278041 459493 278053 459496
rect 278087 459493 278099 459527
rect 278041 459487 278099 459493
rect 287701 459527 287759 459533
rect 287701 459493 287713 459527
rect 287747 459524 287759 459527
rect 296625 459527 296683 459533
rect 296625 459524 296637 459527
rect 287747 459496 296637 459524
rect 287747 459493 287759 459496
rect 287701 459487 287759 459493
rect 296625 459493 296637 459496
rect 296671 459493 296683 459527
rect 296625 459487 296683 459493
rect 306377 459527 306435 459533
rect 306377 459493 306389 459527
rect 306423 459524 306435 459527
rect 315945 459527 316003 459533
rect 315945 459524 315957 459527
rect 306423 459496 315957 459524
rect 306423 459493 306435 459496
rect 306377 459487 306435 459493
rect 315945 459493 315957 459496
rect 315991 459493 316003 459527
rect 315945 459487 316003 459493
rect 6917 459459 6975 459465
rect 6917 459425 6929 459459
rect 6963 459456 6975 459459
rect 16485 459459 16543 459465
rect 16485 459456 16497 459459
rect 6963 459428 16497 459456
rect 6963 459425 6975 459428
rect 6917 459419 6975 459425
rect 16485 459425 16497 459428
rect 16531 459425 16543 459459
rect 16485 459419 16543 459425
rect 26237 459459 26295 459465
rect 26237 459425 26249 459459
rect 26283 459456 26295 459459
rect 35805 459459 35863 459465
rect 35805 459456 35817 459459
rect 26283 459428 35817 459456
rect 26283 459425 26295 459428
rect 26237 459419 26295 459425
rect 35805 459425 35817 459428
rect 35851 459425 35863 459459
rect 35805 459419 35863 459425
rect 45557 459459 45615 459465
rect 45557 459425 45569 459459
rect 45603 459456 45615 459459
rect 55125 459459 55183 459465
rect 55125 459456 55137 459459
rect 45603 459428 55137 459456
rect 45603 459425 45615 459428
rect 45557 459419 45615 459425
rect 55125 459425 55137 459428
rect 55171 459425 55183 459459
rect 55125 459419 55183 459425
rect 64877 459459 64935 459465
rect 64877 459425 64889 459459
rect 64923 459456 64935 459459
rect 74445 459459 74503 459465
rect 74445 459456 74457 459459
rect 64923 459428 74457 459456
rect 64923 459425 64935 459428
rect 64877 459419 64935 459425
rect 74445 459425 74457 459428
rect 74491 459425 74503 459459
rect 74445 459419 74503 459425
rect 84841 459459 84899 459465
rect 84841 459425 84853 459459
rect 84887 459456 84899 459459
rect 94501 459459 94559 459465
rect 94501 459456 94513 459459
rect 84887 459428 94513 459456
rect 84887 459425 84899 459428
rect 84841 459419 84899 459425
rect 94501 459425 94513 459428
rect 94547 459425 94559 459459
rect 94501 459419 94559 459425
rect 104161 459459 104219 459465
rect 104161 459425 104173 459459
rect 104207 459456 104219 459459
rect 113821 459459 113879 459465
rect 113821 459456 113833 459459
rect 104207 459428 113833 459456
rect 104207 459425 104219 459428
rect 104161 459419 104219 459425
rect 113821 459425 113833 459428
rect 113867 459425 113879 459459
rect 113821 459419 113879 459425
rect 123481 459459 123539 459465
rect 123481 459425 123493 459459
rect 123527 459456 123539 459459
rect 133141 459459 133199 459465
rect 133141 459456 133153 459459
rect 123527 459428 133153 459456
rect 123527 459425 123539 459428
rect 123481 459419 123539 459425
rect 133141 459425 133153 459428
rect 133187 459425 133199 459459
rect 133141 459419 133199 459425
rect 142801 459459 142859 459465
rect 142801 459425 142813 459459
rect 142847 459456 142859 459459
rect 152461 459459 152519 459465
rect 152461 459456 152473 459459
rect 142847 459428 152473 459456
rect 142847 459425 142859 459428
rect 142801 459419 142859 459425
rect 152461 459425 152473 459428
rect 152507 459425 152519 459459
rect 152461 459419 152519 459425
rect 162121 459459 162179 459465
rect 162121 459425 162133 459459
rect 162167 459456 162179 459459
rect 171781 459459 171839 459465
rect 171781 459456 171793 459459
rect 162167 459428 171793 459456
rect 162167 459425 162179 459428
rect 162121 459419 162179 459425
rect 171781 459425 171793 459428
rect 171827 459425 171839 459459
rect 171781 459419 171839 459425
rect 181441 459459 181499 459465
rect 181441 459425 181453 459459
rect 181487 459456 181499 459459
rect 191101 459459 191159 459465
rect 191101 459456 191113 459459
rect 181487 459428 191113 459456
rect 181487 459425 181499 459428
rect 181441 459419 181499 459425
rect 191101 459425 191113 459428
rect 191147 459425 191159 459459
rect 191101 459419 191159 459425
rect 200761 459459 200819 459465
rect 200761 459425 200773 459459
rect 200807 459456 200819 459459
rect 210421 459459 210479 459465
rect 210421 459456 210433 459459
rect 200807 459428 210433 459456
rect 200807 459425 200819 459428
rect 200761 459419 200819 459425
rect 210421 459425 210433 459428
rect 210467 459425 210479 459459
rect 210421 459419 210479 459425
rect 220081 459459 220139 459465
rect 220081 459425 220093 459459
rect 220127 459456 220139 459459
rect 225325 459459 225383 459465
rect 225325 459456 225337 459459
rect 220127 459428 225337 459456
rect 220127 459425 220139 459428
rect 220081 459419 220139 459425
rect 225325 459425 225337 459428
rect 225371 459425 225383 459459
rect 238018 459456 238024 459468
rect 237979 459428 238024 459456
rect 225325 459419 225383 459425
rect 238018 459416 238024 459428
rect 238076 459416 238082 459468
rect 240042 459456 240048 459468
rect 240003 459428 240048 459456
rect 240042 459416 240048 459428
rect 240100 459416 240106 459468
rect 243354 459456 243360 459468
rect 243315 459428 243360 459456
rect 243354 459416 243360 459428
rect 243412 459416 243418 459468
rect 246482 459456 246488 459468
rect 246443 459428 246488 459456
rect 246482 459416 246488 459428
rect 246540 459416 246546 459468
rect 249610 459456 249616 459468
rect 249571 459428 249616 459456
rect 249610 459416 249616 459428
rect 249668 459416 249674 459468
rect 254946 459456 254952 459468
rect 254907 459428 254952 459456
rect 254946 459416 254952 459428
rect 255004 459416 255010 459468
rect 257982 459416 257988 459468
rect 258040 459456 258046 459468
rect 349890 459456 349896 459468
rect 258040 459428 349896 459456
rect 258040 459416 258046 459428
rect 349890 459416 349896 459428
rect 349948 459416 349954 459468
rect 3050 459348 3056 459400
rect 3108 459388 3114 459400
rect 321646 459388 321652 459400
rect 3108 459360 321652 459388
rect 3108 459348 3114 459360
rect 321646 459348 321652 459360
rect 321704 459348 321710 459400
rect 329006 459388 329012 459400
rect 327460 459360 329012 459388
rect 4062 459280 4068 459332
rect 4120 459320 4126 459332
rect 325878 459320 325884 459332
rect 4120 459292 325884 459320
rect 4120 459280 4126 459292
rect 325878 459280 325884 459292
rect 325936 459280 325942 459332
rect 16485 459255 16543 459261
rect 16485 459221 16497 459255
rect 16531 459252 16543 459255
rect 16577 459255 16635 459261
rect 16577 459252 16589 459255
rect 16531 459224 16589 459252
rect 16531 459221 16543 459224
rect 16485 459215 16543 459221
rect 16577 459221 16589 459224
rect 16623 459221 16635 459255
rect 16577 459215 16635 459221
rect 35805 459255 35863 459261
rect 35805 459221 35817 459255
rect 35851 459252 35863 459255
rect 35897 459255 35955 459261
rect 35897 459252 35909 459255
rect 35851 459224 35909 459252
rect 35851 459221 35863 459224
rect 35805 459215 35863 459221
rect 35897 459221 35909 459224
rect 35943 459221 35955 459255
rect 35897 459215 35955 459221
rect 55125 459255 55183 459261
rect 55125 459221 55137 459255
rect 55171 459252 55183 459255
rect 55217 459255 55275 459261
rect 55217 459252 55229 459255
rect 55171 459224 55229 459252
rect 55171 459221 55183 459224
rect 55125 459215 55183 459221
rect 55217 459221 55229 459224
rect 55263 459221 55275 459255
rect 55217 459215 55275 459221
rect 74445 459255 74503 459261
rect 74445 459221 74457 459255
rect 74491 459252 74503 459255
rect 74537 459255 74595 459261
rect 74537 459252 74549 459255
rect 74491 459224 74549 459252
rect 74491 459221 74503 459224
rect 74445 459215 74503 459221
rect 74537 459221 74549 459224
rect 74583 459221 74595 459255
rect 74537 459215 74595 459221
rect 234617 459255 234675 459261
rect 234617 459221 234629 459255
rect 234663 459252 234675 459255
rect 247405 459255 247463 459261
rect 247405 459252 247417 459255
rect 234663 459224 247417 459252
rect 234663 459221 234675 459224
rect 234617 459215 234675 459221
rect 247405 459221 247417 459224
rect 247451 459221 247463 459255
rect 247405 459215 247463 459221
rect 258721 459255 258779 459261
rect 258721 459221 258733 459255
rect 258767 459252 258779 459255
rect 268381 459255 268439 459261
rect 268381 459252 268393 459255
rect 258767 459224 268393 459252
rect 258767 459221 258779 459224
rect 258721 459215 258779 459221
rect 268381 459221 268393 459224
rect 268427 459221 268439 459255
rect 268381 459215 268439 459221
rect 278041 459255 278099 459261
rect 278041 459221 278053 459255
rect 278087 459252 278099 459255
rect 287701 459255 287759 459261
rect 287701 459252 287713 459255
rect 278087 459224 287713 459252
rect 278087 459221 278099 459224
rect 278041 459215 278099 459221
rect 287701 459221 287713 459224
rect 287747 459221 287759 459255
rect 287701 459215 287759 459221
rect 296625 459255 296683 459261
rect 296625 459221 296637 459255
rect 296671 459252 296683 459255
rect 306377 459255 306435 459261
rect 306377 459252 306389 459255
rect 296671 459224 306389 459252
rect 296671 459221 296683 459224
rect 296625 459215 296683 459221
rect 306377 459221 306389 459224
rect 306423 459221 306435 459255
rect 306377 459215 306435 459221
rect 315945 459255 316003 459261
rect 315945 459221 315957 459255
rect 315991 459252 316003 459255
rect 327460 459252 327488 459360
rect 329006 459348 329012 459360
rect 329064 459348 329070 459400
rect 327902 459280 327908 459332
rect 327960 459280 327966 459332
rect 331214 459320 331220 459332
rect 331175 459292 331220 459320
rect 331214 459280 331220 459292
rect 331272 459280 331278 459332
rect 332134 459320 332140 459332
rect 332095 459292 332140 459320
rect 332134 459280 332140 459292
rect 332192 459280 332198 459332
rect 334158 459320 334164 459332
rect 334119 459292 334164 459320
rect 334158 459280 334164 459292
rect 334216 459280 334222 459332
rect 335354 459280 335360 459332
rect 335412 459320 335418 459332
rect 337286 459320 337292 459332
rect 335412 459292 335457 459320
rect 337247 459292 337292 459320
rect 335412 459280 335418 459292
rect 337286 459280 337292 459292
rect 337344 459280 337350 459332
rect 338390 459320 338396 459332
rect 338351 459292 338396 459320
rect 338390 459280 338396 459292
rect 338448 459280 338454 459332
rect 340690 459320 340696 459332
rect 340651 459292 340696 459320
rect 340690 459280 340696 459292
rect 340748 459280 340754 459332
rect 341518 459320 341524 459332
rect 341479 459292 341524 459320
rect 341518 459280 341524 459292
rect 341576 459280 341582 459332
rect 315991 459224 327488 459252
rect 315991 459221 316003 459224
rect 315945 459215 316003 459221
rect 3970 459144 3976 459196
rect 4028 459184 4034 459196
rect 327920 459184 327948 459280
rect 4028 459156 327948 459184
rect 4028 459144 4034 459156
rect 5350 459076 5356 459128
rect 5408 459116 5414 459128
rect 6917 459119 6975 459125
rect 6917 459116 6929 459119
rect 5408 459088 6929 459116
rect 5408 459076 5414 459088
rect 6917 459085 6929 459088
rect 6963 459085 6975 459119
rect 6917 459079 6975 459085
rect 16577 459119 16635 459125
rect 16577 459085 16589 459119
rect 16623 459116 16635 459119
rect 26237 459119 26295 459125
rect 26237 459116 26249 459119
rect 16623 459088 26249 459116
rect 16623 459085 16635 459088
rect 16577 459079 16635 459085
rect 26237 459085 26249 459088
rect 26283 459085 26295 459119
rect 26237 459079 26295 459085
rect 35897 459119 35955 459125
rect 35897 459085 35909 459119
rect 35943 459116 35955 459119
rect 45557 459119 45615 459125
rect 45557 459116 45569 459119
rect 35943 459088 45569 459116
rect 35943 459085 35955 459088
rect 35897 459079 35955 459085
rect 45557 459085 45569 459088
rect 45603 459085 45615 459119
rect 45557 459079 45615 459085
rect 55217 459119 55275 459125
rect 55217 459085 55229 459119
rect 55263 459116 55275 459119
rect 64877 459119 64935 459125
rect 64877 459116 64889 459119
rect 55263 459088 64889 459116
rect 55263 459085 55275 459088
rect 55217 459079 55275 459085
rect 64877 459085 64889 459088
rect 64923 459085 64935 459119
rect 64877 459079 64935 459085
rect 74537 459119 74595 459125
rect 74537 459085 74549 459119
rect 74583 459116 74595 459119
rect 84841 459119 84899 459125
rect 84841 459116 84853 459119
rect 74583 459088 84853 459116
rect 74583 459085 74595 459088
rect 74537 459079 74595 459085
rect 84841 459085 84853 459088
rect 84887 459085 84899 459119
rect 84841 459079 84899 459085
rect 94501 459119 94559 459125
rect 94501 459085 94513 459119
rect 94547 459116 94559 459119
rect 104161 459119 104219 459125
rect 104161 459116 104173 459119
rect 94547 459088 104173 459116
rect 94547 459085 94559 459088
rect 94501 459079 94559 459085
rect 104161 459085 104173 459088
rect 104207 459085 104219 459119
rect 104161 459079 104219 459085
rect 113821 459119 113879 459125
rect 113821 459085 113833 459119
rect 113867 459116 113879 459119
rect 123481 459119 123539 459125
rect 123481 459116 123493 459119
rect 113867 459088 123493 459116
rect 113867 459085 113879 459088
rect 113821 459079 113879 459085
rect 123481 459085 123493 459088
rect 123527 459085 123539 459119
rect 123481 459079 123539 459085
rect 133141 459119 133199 459125
rect 133141 459085 133153 459119
rect 133187 459116 133199 459119
rect 142801 459119 142859 459125
rect 142801 459116 142813 459119
rect 133187 459088 142813 459116
rect 133187 459085 133199 459088
rect 133141 459079 133199 459085
rect 142801 459085 142813 459088
rect 142847 459085 142859 459119
rect 142801 459079 142859 459085
rect 152461 459119 152519 459125
rect 152461 459085 152473 459119
rect 152507 459116 152519 459119
rect 162121 459119 162179 459125
rect 162121 459116 162133 459119
rect 152507 459088 162133 459116
rect 152507 459085 152519 459088
rect 152461 459079 152519 459085
rect 162121 459085 162133 459088
rect 162167 459085 162179 459119
rect 162121 459079 162179 459085
rect 171781 459119 171839 459125
rect 171781 459085 171793 459119
rect 171827 459116 171839 459119
rect 181441 459119 181499 459125
rect 181441 459116 181453 459119
rect 171827 459088 181453 459116
rect 171827 459085 171839 459088
rect 171781 459079 171839 459085
rect 181441 459085 181453 459088
rect 181487 459085 181499 459119
rect 181441 459079 181499 459085
rect 191101 459119 191159 459125
rect 191101 459085 191113 459119
rect 191147 459116 191159 459119
rect 200761 459119 200819 459125
rect 200761 459116 200773 459119
rect 191147 459088 200773 459116
rect 191147 459085 191159 459088
rect 191101 459079 191159 459085
rect 200761 459085 200773 459088
rect 200807 459085 200819 459119
rect 200761 459079 200819 459085
rect 210421 459119 210479 459125
rect 210421 459085 210433 459119
rect 210467 459116 210479 459119
rect 220081 459119 220139 459125
rect 220081 459116 220093 459119
rect 210467 459088 220093 459116
rect 210467 459085 210479 459088
rect 210421 459079 210479 459085
rect 220081 459085 220093 459088
rect 220127 459085 220139 459119
rect 220081 459079 220139 459085
rect 225325 459119 225383 459125
rect 225325 459085 225337 459119
rect 225371 459116 225383 459119
rect 234617 459119 234675 459125
rect 234617 459116 234629 459119
rect 225371 459088 234629 459116
rect 225371 459085 225383 459088
rect 225325 459079 225383 459085
rect 234617 459085 234629 459088
rect 234663 459085 234675 459119
rect 234617 459079 234675 459085
rect 254949 459119 255007 459125
rect 254949 459085 254961 459119
rect 254995 459116 255007 459119
rect 579890 459116 579896 459128
rect 254995 459088 579896 459116
rect 254995 459085 255007 459088
rect 254949 459079 255007 459085
rect 579890 459076 579896 459088
rect 579948 459076 579954 459128
rect 5166 459008 5172 459060
rect 5224 459048 5230 459060
rect 332137 459051 332195 459057
rect 332137 459048 332149 459051
rect 5224 459020 332149 459048
rect 5224 459008 5230 459020
rect 332137 459017 332149 459020
rect 332183 459017 332195 459051
rect 332137 459011 332195 459017
rect 3878 458940 3884 458992
rect 3936 458980 3942 458992
rect 331217 458983 331275 458989
rect 331217 458980 331229 458983
rect 3936 458952 331229 458980
rect 3936 458940 3942 458952
rect 331217 458949 331229 458952
rect 331263 458949 331275 458983
rect 331217 458943 331275 458949
rect 3786 458872 3792 458924
rect 3844 458912 3850 458924
rect 334161 458915 334219 458921
rect 334161 458912 334173 458915
rect 3844 458884 334173 458912
rect 3844 458872 3850 458884
rect 334161 458881 334173 458884
rect 334207 458881 334219 458915
rect 334161 458875 334219 458881
rect 249613 458847 249671 458853
rect 249613 458813 249625 458847
rect 249659 458844 249671 458847
rect 580074 458844 580080 458856
rect 249659 458816 580080 458844
rect 249659 458813 249671 458816
rect 249613 458807 249671 458813
rect 580074 458804 580080 458816
rect 580132 458804 580138 458856
rect 4982 458736 4988 458788
rect 5040 458776 5046 458788
rect 335357 458779 335415 458785
rect 335357 458776 335369 458779
rect 5040 458748 335369 458776
rect 5040 458736 5046 458748
rect 335357 458745 335369 458748
rect 335403 458745 335415 458779
rect 335357 458739 335415 458745
rect 3694 458668 3700 458720
rect 3752 458708 3758 458720
rect 337289 458711 337347 458717
rect 337289 458708 337301 458711
rect 3752 458680 337301 458708
rect 3752 458668 3758 458680
rect 337289 458677 337301 458680
rect 337335 458677 337347 458711
rect 337289 458671 337347 458677
rect 4798 458600 4804 458652
rect 4856 458640 4862 458652
rect 338393 458643 338451 458649
rect 338393 458640 338405 458643
rect 4856 458612 338405 458640
rect 4856 458600 4862 458612
rect 338393 458609 338405 458612
rect 338439 458609 338451 458643
rect 338393 458603 338451 458609
rect 246485 458575 246543 458581
rect 246485 458541 246497 458575
rect 246531 458572 246543 458575
rect 580902 458572 580908 458584
rect 246531 458544 580908 458572
rect 246531 458541 246543 458544
rect 246485 458535 246543 458541
rect 580902 458532 580908 458544
rect 580960 458532 580966 458584
rect 243357 458507 243415 458513
rect 243357 458473 243369 458507
rect 243403 458504 243415 458507
rect 580718 458504 580724 458516
rect 243403 458476 580724 458504
rect 243403 458473 243415 458476
rect 243357 458467 243415 458473
rect 580718 458464 580724 458476
rect 580776 458464 580782 458516
rect 3602 458396 3608 458448
rect 3660 458436 3666 458448
rect 340693 458439 340751 458445
rect 340693 458436 340705 458439
rect 3660 458408 340705 458436
rect 3660 458396 3666 458408
rect 340693 458405 340705 458408
rect 340739 458405 340751 458439
rect 340693 458399 340751 458405
rect 3510 458328 3516 458380
rect 3568 458368 3574 458380
rect 341521 458371 341579 458377
rect 341521 458368 341533 458371
rect 3568 458340 341533 458368
rect 3568 458328 3574 458340
rect 341521 458337 341533 458340
rect 341567 458337 341579 458371
rect 341521 458331 341579 458337
rect 240045 458303 240103 458309
rect 240045 458269 240057 458303
rect 240091 458300 240103 458303
rect 580534 458300 580540 458312
rect 240091 458272 580540 458300
rect 240091 458269 240103 458272
rect 240045 458263 240103 458269
rect 580534 458260 580540 458272
rect 580592 458260 580598 458312
rect 238021 458235 238079 458241
rect 238021 458201 238033 458235
rect 238067 458232 238079 458235
rect 580442 458232 580448 458244
rect 238067 458204 580448 458232
rect 238067 458201 238079 458204
rect 238021 458195 238079 458201
rect 580442 458192 580448 458204
rect 580500 458192 580506 458244
rect 579706 451596 579712 451648
rect 579764 451636 579770 451648
rect 580166 451636 580172 451648
rect 579764 451608 580172 451636
rect 579764 451596 579770 451608
rect 580166 451596 580172 451608
rect 580224 451596 580230 451648
rect 2774 437996 2780 438048
rect 2832 438036 2838 438048
rect 4614 438036 4620 438048
rect 2832 438008 4620 438036
rect 2832 437996 2838 438008
rect 4614 437996 4620 438008
rect 4672 437996 4678 438048
rect 349890 405628 349896 405680
rect 349948 405668 349954 405680
rect 579798 405668 579804 405680
rect 349948 405640 579804 405668
rect 349948 405628 349954 405640
rect 579798 405628 579804 405640
rect 579856 405628 579862 405680
rect 281718 340144 281724 340196
rect 281776 340184 281782 340196
rect 282454 340184 282460 340196
rect 281776 340156 282460 340184
rect 281776 340144 281782 340156
rect 282454 340144 282460 340156
rect 282512 340144 282518 340196
rect 299566 340144 299572 340196
rect 299624 340184 299630 340196
rect 300578 340184 300584 340196
rect 299624 340156 300584 340184
rect 299624 340144 299630 340156
rect 300578 340144 300584 340156
rect 300636 340144 300642 340196
rect 317877 340187 317935 340193
rect 317877 340153 317889 340187
rect 317923 340184 317935 340187
rect 317966 340184 317972 340196
rect 317923 340156 317972 340184
rect 317923 340153 317935 340156
rect 317877 340147 317935 340153
rect 317966 340144 317972 340156
rect 318024 340144 318030 340196
rect 262582 339056 262588 339108
rect 262640 339096 262646 339108
rect 263042 339096 263048 339108
rect 262640 339068 263048 339096
rect 262640 339056 262646 339068
rect 263042 339056 263048 339068
rect 263100 339056 263106 339108
rect 270678 339056 270684 339108
rect 270736 339096 270742 339108
rect 271138 339096 271144 339108
rect 270736 339068 271144 339096
rect 270736 339056 270742 339068
rect 271138 339056 271144 339068
rect 271196 339056 271202 339108
rect 302970 339056 302976 339108
rect 303028 339096 303034 339108
rect 303338 339096 303344 339108
rect 303028 339068 303344 339096
rect 303028 339056 303034 339068
rect 303338 339056 303344 339068
rect 303396 339056 303402 339108
rect 243354 338920 243360 338972
rect 243412 338960 243418 338972
rect 243722 338960 243728 338972
rect 243412 338932 243728 338960
rect 243412 338920 243418 338932
rect 243722 338920 243728 338932
rect 243780 338920 243786 338972
rect 267734 338920 267740 338972
rect 267792 338960 267798 338972
rect 268194 338960 268200 338972
rect 267792 338932 268200 338960
rect 267792 338920 267798 338932
rect 268194 338920 268200 338932
rect 268252 338920 268258 338972
rect 309134 338920 309140 338972
rect 309192 338960 309198 338972
rect 309502 338960 309508 338972
rect 309192 338932 309508 338960
rect 309192 338920 309198 338932
rect 309502 338920 309508 338932
rect 309560 338920 309566 338972
rect 316494 338920 316500 338972
rect 316552 338960 316558 338972
rect 316862 338960 316868 338972
rect 316552 338932 316868 338960
rect 316552 338920 316558 338932
rect 316862 338920 316868 338932
rect 316920 338920 316926 338972
rect 258718 338852 258724 338904
rect 258776 338892 258782 338904
rect 259086 338892 259092 338904
rect 258776 338864 259092 338892
rect 258776 338852 258782 338864
rect 259086 338852 259092 338864
rect 259144 338852 259150 338904
rect 232866 338784 232872 338836
rect 232924 338824 232930 338836
rect 233142 338824 233148 338836
rect 232924 338796 233148 338824
rect 232924 338784 232930 338796
rect 233142 338784 233148 338796
rect 233200 338784 233206 338836
rect 241698 338784 241704 338836
rect 241756 338824 241762 338836
rect 242066 338824 242072 338836
rect 241756 338796 242072 338824
rect 241756 338784 241762 338796
rect 242066 338784 242072 338796
rect 242124 338784 242130 338836
rect 231854 338648 231860 338700
rect 231912 338688 231918 338700
rect 232130 338688 232136 338700
rect 231912 338660 232136 338688
rect 231912 338648 231918 338660
rect 232130 338648 232136 338660
rect 232188 338648 232194 338700
rect 238018 338648 238024 338700
rect 238076 338688 238082 338700
rect 238294 338688 238300 338700
rect 238076 338660 238300 338688
rect 238076 338648 238082 338660
rect 238294 338648 238300 338660
rect 238352 338648 238358 338700
rect 259454 338648 259460 338700
rect 259512 338688 259518 338700
rect 259822 338688 259828 338700
rect 259512 338660 259828 338688
rect 259512 338648 259518 338660
rect 259822 338648 259828 338660
rect 259880 338648 259886 338700
rect 343726 338648 343732 338700
rect 343784 338688 343790 338700
rect 344094 338688 344100 338700
rect 343784 338660 344100 338688
rect 343784 338648 343790 338660
rect 344094 338648 344100 338660
rect 344152 338648 344158 338700
rect 242986 338512 242992 338564
rect 243044 338552 243050 338564
rect 243262 338552 243268 338564
rect 243044 338524 243268 338552
rect 243044 338512 243050 338524
rect 243262 338512 243268 338524
rect 243320 338512 243326 338564
rect 334158 338512 334164 338564
rect 334216 338552 334222 338564
rect 334526 338552 334532 338564
rect 334216 338524 334532 338552
rect 334216 338512 334222 338524
rect 334526 338512 334532 338524
rect 334584 338512 334590 338564
rect 272150 338376 272156 338428
rect 272208 338416 272214 338428
rect 272610 338416 272616 338428
rect 272208 338388 272616 338416
rect 272208 338376 272214 338388
rect 272610 338376 272616 338388
rect 272668 338376 272674 338428
rect 280246 338376 280252 338428
rect 280304 338416 280310 338428
rect 280614 338416 280620 338428
rect 280304 338388 280620 338416
rect 280304 338376 280310 338388
rect 280614 338376 280620 338388
rect 280672 338376 280678 338428
rect 287238 338376 287244 338428
rect 287296 338416 287302 338428
rect 287698 338416 287704 338428
rect 287296 338388 287704 338416
rect 287296 338376 287302 338388
rect 287698 338376 287704 338388
rect 287756 338376 287762 338428
rect 289998 338376 290004 338428
rect 290056 338416 290062 338428
rect 290274 338416 290280 338428
rect 290056 338388 290280 338416
rect 290056 338376 290062 338388
rect 290274 338376 290280 338388
rect 290332 338376 290338 338428
rect 341058 338376 341064 338428
rect 341116 338416 341122 338428
rect 341334 338416 341340 338428
rect 341116 338388 341340 338416
rect 341116 338376 341122 338388
rect 341334 338376 341340 338388
rect 341392 338376 341398 338428
rect 309870 338104 309876 338156
rect 309928 338144 309934 338156
rect 310054 338144 310060 338156
rect 309928 338116 310060 338144
rect 309928 338104 309934 338116
rect 310054 338104 310060 338116
rect 310112 338104 310118 338156
rect 317874 338144 317880 338156
rect 317835 338116 317880 338144
rect 317874 338104 317880 338116
rect 317932 338104 317938 338156
rect 319530 338104 319536 338156
rect 319588 338144 319594 338156
rect 320082 338144 320088 338156
rect 319588 338116 320088 338144
rect 319588 338104 319594 338116
rect 320082 338104 320088 338116
rect 320140 338104 320146 338156
rect 86862 338036 86868 338088
rect 86920 338076 86926 338088
rect 341610 338076 341616 338088
rect 86920 338048 341616 338076
rect 86920 338036 86926 338048
rect 341610 338036 341616 338048
rect 341668 338036 341674 338088
rect 93762 337968 93768 338020
rect 93820 338008 93826 338020
rect 343082 338008 343088 338020
rect 93820 337980 343088 338008
rect 93820 337968 93826 337980
rect 343082 337968 343088 337980
rect 343140 337968 343146 338020
rect 82722 337900 82728 337952
rect 82780 337940 82786 337952
rect 340874 337940 340880 337952
rect 82780 337912 340880 337940
rect 82780 337900 82786 337912
rect 340874 337900 340880 337912
rect 340932 337900 340938 337952
rect 75822 337832 75828 337884
rect 75880 337872 75886 337884
rect 339402 337872 339408 337884
rect 75880 337844 339408 337872
rect 75880 337832 75886 337844
rect 339402 337832 339408 337844
rect 339460 337832 339466 337884
rect 62022 337764 62028 337816
rect 62080 337804 62086 337816
rect 336458 337804 336464 337816
rect 62080 337776 336464 337804
rect 62080 337764 62086 337776
rect 336458 337764 336464 337776
rect 336516 337764 336522 337816
rect 68922 337696 68928 337748
rect 68980 337736 68986 337748
rect 337930 337736 337936 337748
rect 68980 337708 337936 337736
rect 68980 337696 68986 337708
rect 337930 337696 337936 337708
rect 337988 337696 337994 337748
rect 57882 337628 57888 337680
rect 57940 337668 57946 337680
rect 335722 337668 335728 337680
rect 57940 337640 335728 337668
rect 57940 337628 57946 337640
rect 335722 337628 335728 337640
rect 335780 337628 335786 337680
rect 44082 337560 44088 337612
rect 44140 337600 44146 337612
rect 44140 337572 331076 337600
rect 44140 337560 44146 337572
rect 55122 337492 55128 337544
rect 55180 337532 55186 337544
rect 326433 337535 326491 337541
rect 55180 337504 326384 337532
rect 55180 337492 55186 337504
rect 42702 337424 42708 337476
rect 42760 337464 42766 337476
rect 42760 337436 322980 337464
rect 42760 337424 42766 337436
rect 35802 337356 35808 337408
rect 35860 337396 35866 337408
rect 322014 337396 322020 337408
rect 35860 337368 322020 337396
rect 35860 337356 35866 337368
rect 322014 337356 322020 337368
rect 322072 337356 322078 337408
rect 322198 337356 322204 337408
rect 322256 337396 322262 337408
rect 322750 337396 322756 337408
rect 322256 337368 322756 337396
rect 322256 337356 322262 337368
rect 322750 337356 322756 337368
rect 322808 337356 322814 337408
rect 322952 337396 322980 337436
rect 323118 337424 323124 337476
rect 323176 337464 323182 337476
rect 323762 337464 323768 337476
rect 323176 337436 323768 337464
rect 323176 337424 323182 337436
rect 323762 337424 323768 337436
rect 323820 337424 323826 337476
rect 323946 337424 323952 337476
rect 324004 337464 324010 337476
rect 326249 337467 326307 337473
rect 326249 337464 326261 337467
rect 324004 337436 326261 337464
rect 324004 337424 324010 337436
rect 326249 337433 326261 337436
rect 326295 337433 326307 337467
rect 326356 337464 326384 337504
rect 326433 337501 326445 337535
rect 326479 337532 326491 337535
rect 330938 337532 330944 337544
rect 326479 337504 330944 337532
rect 326479 337501 326491 337504
rect 326433 337495 326491 337501
rect 330938 337492 330944 337504
rect 330996 337492 331002 337544
rect 331048 337532 331076 337572
rect 332778 337532 332784 337544
rect 331048 337504 332784 337532
rect 332778 337492 332784 337504
rect 332836 337492 332842 337544
rect 331125 337467 331183 337473
rect 331125 337464 331137 337467
rect 326356 337436 331137 337464
rect 326249 337427 326307 337433
rect 331125 337433 331137 337436
rect 331171 337433 331183 337467
rect 331125 337427 331183 337433
rect 331217 337467 331275 337473
rect 331217 337433 331229 337467
rect 331263 337464 331275 337467
rect 334986 337464 334992 337476
rect 331263 337436 334992 337464
rect 331263 337433 331275 337436
rect 331217 337427 331275 337433
rect 334986 337424 334992 337436
rect 335044 337424 335050 337476
rect 332594 337396 332600 337408
rect 322952 337368 332600 337396
rect 332594 337356 332600 337368
rect 332652 337356 332658 337408
rect 100662 337288 100668 337340
rect 100720 337328 100726 337340
rect 344554 337328 344560 337340
rect 100720 337300 344560 337328
rect 100720 337288 100726 337300
rect 344554 337288 344560 337300
rect 344612 337288 344618 337340
rect 107470 337220 107476 337272
rect 107528 337260 107534 337272
rect 346026 337260 346032 337272
rect 107528 337232 346032 337260
rect 107528 337220 107534 337232
rect 346026 337220 346032 337232
rect 346084 337220 346090 337272
rect 115842 337152 115848 337204
rect 115900 337192 115906 337204
rect 347498 337192 347504 337204
rect 115900 337164 347504 337192
rect 115900 337152 115906 337164
rect 347498 337152 347504 337164
rect 347556 337152 347562 337204
rect 122742 337084 122748 337136
rect 122800 337124 122806 337136
rect 348970 337124 348976 337136
rect 122800 337096 348976 337124
rect 122800 337084 122806 337096
rect 348970 337084 348976 337096
rect 349028 337084 349034 337136
rect 173158 337016 173164 337068
rect 173216 337056 173222 337068
rect 345750 337056 345756 337068
rect 173216 337028 345756 337056
rect 173216 337016 173222 337028
rect 345750 337016 345756 337028
rect 345808 337016 345814 337068
rect 182818 336948 182824 337000
rect 182876 336988 182882 337000
rect 347222 336988 347228 337000
rect 182876 336960 347228 336988
rect 182876 336948 182882 336960
rect 347222 336948 347228 336960
rect 347280 336948 347286 337000
rect 186958 336880 186964 336932
rect 187016 336920 187022 336932
rect 348694 336920 348700 336932
rect 187016 336892 348700 336920
rect 187016 336880 187022 336892
rect 348694 336880 348700 336892
rect 348752 336880 348758 336932
rect 191098 336812 191104 336864
rect 191156 336852 191162 336864
rect 349430 336852 349436 336864
rect 191156 336824 349436 336852
rect 191156 336812 191162 336824
rect 349430 336812 349436 336824
rect 349488 336812 349494 336864
rect 195238 336744 195244 336796
rect 195296 336784 195302 336796
rect 349706 336784 349712 336796
rect 195296 336756 349712 336784
rect 195296 336744 195302 336756
rect 349706 336744 349712 336756
rect 349764 336744 349770 336796
rect 107470 336716 107476 336728
rect 107431 336688 107476 336716
rect 107470 336676 107476 336688
rect 107528 336676 107534 336728
rect 271966 336676 271972 336728
rect 272024 336716 272030 336728
rect 272150 336716 272156 336728
rect 272024 336688 272156 336716
rect 272024 336676 272030 336688
rect 272150 336676 272156 336688
rect 272208 336676 272214 336728
rect 279510 336716 279516 336728
rect 279471 336688 279516 336716
rect 279510 336676 279516 336688
rect 279568 336676 279574 336728
rect 305362 336676 305368 336728
rect 305420 336716 305426 336728
rect 305546 336716 305552 336728
rect 305420 336688 305552 336716
rect 305420 336676 305426 336688
rect 305546 336676 305552 336688
rect 305604 336676 305610 336728
rect 331125 336719 331183 336725
rect 331125 336685 331137 336719
rect 331171 336716 331183 336719
rect 331217 336719 331275 336725
rect 331217 336716 331229 336719
rect 331171 336688 331229 336716
rect 331171 336685 331183 336688
rect 331125 336679 331183 336685
rect 331217 336685 331229 336688
rect 331263 336685 331275 336719
rect 331217 336679 331275 336685
rect 291378 336608 291384 336660
rect 291436 336648 291442 336660
rect 291746 336648 291752 336660
rect 291436 336620 291752 336648
rect 291436 336608 291442 336620
rect 291746 336608 291752 336620
rect 291804 336608 291810 336660
rect 313366 335996 313372 336048
rect 313424 336036 313430 336048
rect 313642 336036 313648 336048
rect 313424 336008 313648 336036
rect 313424 335996 313430 336008
rect 313642 335996 313648 336008
rect 313700 335996 313706 336048
rect 313550 335928 313556 335980
rect 313608 335928 313614 335980
rect 320174 335928 320180 335980
rect 320232 335968 320238 335980
rect 320818 335968 320824 335980
rect 320232 335940 320824 335968
rect 320232 335928 320238 335940
rect 320818 335928 320824 335940
rect 320876 335928 320882 335980
rect 235994 335860 236000 335912
rect 236052 335900 236058 335912
rect 236454 335900 236460 335912
rect 236052 335872 236460 335900
rect 236052 335860 236058 335872
rect 236454 335860 236460 335872
rect 236512 335860 236518 335912
rect 236178 335792 236184 335844
rect 236236 335832 236242 335844
rect 236638 335832 236644 335844
rect 236236 335804 236644 335832
rect 236236 335792 236242 335804
rect 236638 335792 236644 335804
rect 236696 335792 236702 335844
rect 245746 335792 245752 335844
rect 245804 335832 245810 335844
rect 245930 335832 245936 335844
rect 245804 335804 245936 335832
rect 245804 335792 245810 335804
rect 245930 335792 245936 335804
rect 245988 335792 245994 335844
rect 261294 335792 261300 335844
rect 261352 335792 261358 335844
rect 269206 335792 269212 335844
rect 269264 335832 269270 335844
rect 270218 335832 270224 335844
rect 269264 335804 270224 335832
rect 269264 335792 269270 335804
rect 270218 335792 270224 335804
rect 270276 335792 270282 335844
rect 273438 335792 273444 335844
rect 273496 335832 273502 335844
rect 273622 335832 273628 335844
rect 273496 335804 273628 335832
rect 273496 335792 273502 335804
rect 273622 335792 273628 335804
rect 273680 335792 273686 335844
rect 299658 335792 299664 335844
rect 299716 335832 299722 335844
rect 299842 335832 299848 335844
rect 299716 335804 299848 335832
rect 299716 335792 299722 335804
rect 299842 335792 299848 335804
rect 299900 335792 299906 335844
rect 311986 335792 311992 335844
rect 312044 335832 312050 335844
rect 312538 335832 312544 335844
rect 312044 335804 312544 335832
rect 312044 335792 312050 335804
rect 312538 335792 312544 335804
rect 312596 335792 312602 335844
rect 232133 335767 232191 335773
rect 232133 335733 232145 335767
rect 232179 335764 232191 335767
rect 232222 335764 232228 335776
rect 232179 335736 232228 335764
rect 232179 335733 232191 335736
rect 232133 335727 232191 335733
rect 232222 335724 232228 335736
rect 232280 335724 232286 335776
rect 261312 335708 261340 335792
rect 313568 335776 313596 335928
rect 317690 335792 317696 335844
rect 317748 335832 317754 335844
rect 317966 335832 317972 335844
rect 317748 335804 317972 335832
rect 317748 335792 317754 335804
rect 317966 335792 317972 335804
rect 318024 335792 318030 335844
rect 284478 335724 284484 335776
rect 284536 335764 284542 335776
rect 284662 335764 284668 335776
rect 284536 335736 284668 335764
rect 284536 335724 284542 335736
rect 284662 335724 284668 335736
rect 284720 335724 284726 335776
rect 291286 335724 291292 335776
rect 291344 335764 291350 335776
rect 292298 335764 292304 335776
rect 291344 335736 292304 335764
rect 291344 335724 291350 335736
rect 292298 335724 292304 335736
rect 292356 335724 292362 335776
rect 303798 335724 303804 335776
rect 303856 335764 303862 335776
rect 303982 335764 303988 335776
rect 303856 335736 303988 335764
rect 303856 335724 303862 335736
rect 303982 335724 303988 335736
rect 304040 335724 304046 335776
rect 313550 335724 313556 335776
rect 313608 335724 313614 335776
rect 328546 335724 328552 335776
rect 328604 335764 328610 335776
rect 328822 335764 328828 335776
rect 328604 335736 328828 335764
rect 328604 335724 328610 335736
rect 328822 335724 328828 335736
rect 328880 335724 328886 335776
rect 233326 335656 233332 335708
rect 233384 335696 233390 335708
rect 234246 335696 234252 335708
rect 233384 335668 234252 335696
rect 233384 335656 233390 335668
rect 234246 335656 234252 335668
rect 234304 335656 234310 335708
rect 237374 335656 237380 335708
rect 237432 335696 237438 335708
rect 238386 335696 238392 335708
rect 237432 335668 238392 335696
rect 237432 335656 237438 335668
rect 238386 335656 238392 335668
rect 238444 335656 238450 335708
rect 247034 335656 247040 335708
rect 247092 335696 247098 335708
rect 248138 335696 248144 335708
rect 247092 335668 248144 335696
rect 247092 335656 247098 335668
rect 248138 335656 248144 335668
rect 248196 335656 248202 335708
rect 248414 335656 248420 335708
rect 248472 335696 248478 335708
rect 248874 335696 248880 335708
rect 248472 335668 248880 335696
rect 248472 335656 248478 335668
rect 248874 335656 248880 335668
rect 248932 335656 248938 335708
rect 249886 335656 249892 335708
rect 249944 335696 249950 335708
rect 250346 335696 250352 335708
rect 249944 335668 250352 335696
rect 249944 335656 249950 335668
rect 250346 335656 250352 335668
rect 250404 335656 250410 335708
rect 251358 335656 251364 335708
rect 251416 335696 251422 335708
rect 251818 335696 251824 335708
rect 251416 335668 251824 335696
rect 251416 335656 251422 335668
rect 251818 335656 251824 335668
rect 251876 335656 251882 335708
rect 252646 335656 252652 335708
rect 252704 335696 252710 335708
rect 253290 335696 253296 335708
rect 252704 335668 253296 335696
rect 252704 335656 252710 335668
rect 253290 335656 253296 335668
rect 253348 335656 253354 335708
rect 254302 335656 254308 335708
rect 254360 335696 254366 335708
rect 254486 335696 254492 335708
rect 254360 335668 254492 335696
rect 254360 335656 254366 335668
rect 254486 335656 254492 335668
rect 254544 335656 254550 335708
rect 255498 335656 255504 335708
rect 255556 335696 255562 335708
rect 256050 335696 256056 335708
rect 255556 335668 256056 335696
rect 255556 335656 255562 335668
rect 256050 335656 256056 335668
rect 256108 335656 256114 335708
rect 261294 335656 261300 335708
rect 261352 335656 261358 335708
rect 262214 335656 262220 335708
rect 262272 335696 262278 335708
rect 263318 335696 263324 335708
rect 262272 335668 263324 335696
rect 262272 335656 262278 335668
rect 263318 335656 263324 335668
rect 263376 335656 263382 335708
rect 266630 335656 266636 335708
rect 266688 335696 266694 335708
rect 267550 335696 267556 335708
rect 266688 335668 267556 335696
rect 266688 335656 266694 335668
rect 267550 335656 267556 335668
rect 267608 335656 267614 335708
rect 267826 335656 267832 335708
rect 267884 335696 267890 335708
rect 268746 335696 268752 335708
rect 267884 335668 268752 335696
rect 267884 335656 267890 335668
rect 268746 335656 268752 335668
rect 268804 335656 268810 335708
rect 269298 335656 269304 335708
rect 269356 335696 269362 335708
rect 270218 335696 270224 335708
rect 269356 335668 270224 335696
rect 269356 335656 269362 335668
rect 270218 335656 270224 335668
rect 270276 335656 270282 335708
rect 276198 335656 276204 335708
rect 276256 335696 276262 335708
rect 277302 335696 277308 335708
rect 276256 335668 277308 335696
rect 276256 335656 276262 335668
rect 277302 335656 277308 335668
rect 277360 335656 277366 335708
rect 277394 335656 277400 335708
rect 277452 335696 277458 335708
rect 278222 335696 278228 335708
rect 277452 335668 278228 335696
rect 277452 335656 277458 335668
rect 278222 335656 278228 335668
rect 278280 335656 278286 335708
rect 280154 335656 280160 335708
rect 280212 335696 280218 335708
rect 281258 335696 281264 335708
rect 280212 335668 281264 335696
rect 280212 335656 280218 335668
rect 281258 335656 281264 335668
rect 281316 335656 281322 335708
rect 281534 335656 281540 335708
rect 281592 335696 281598 335708
rect 282730 335696 282736 335708
rect 281592 335668 282736 335696
rect 281592 335656 281598 335668
rect 282730 335656 282736 335668
rect 282788 335656 282794 335708
rect 284386 335656 284392 335708
rect 284444 335696 284450 335708
rect 284938 335696 284944 335708
rect 284444 335668 284944 335696
rect 284444 335656 284450 335668
rect 284938 335656 284944 335668
rect 284996 335656 285002 335708
rect 286042 335656 286048 335708
rect 286100 335696 286106 335708
rect 286778 335696 286784 335708
rect 286100 335668 286784 335696
rect 286100 335656 286106 335668
rect 286778 335656 286784 335668
rect 286836 335656 286842 335708
rect 289906 335656 289912 335708
rect 289964 335696 289970 335708
rect 290734 335696 290740 335708
rect 289964 335668 290740 335696
rect 289964 335656 289970 335668
rect 290734 335656 290740 335668
rect 290792 335656 290798 335708
rect 291562 335656 291568 335708
rect 291620 335696 291626 335708
rect 292022 335696 292028 335708
rect 291620 335668 292028 335696
rect 291620 335656 291626 335668
rect 292022 335656 292028 335668
rect 292080 335656 292086 335708
rect 293034 335656 293040 335708
rect 293092 335696 293098 335708
rect 293678 335696 293684 335708
rect 293092 335668 293684 335696
rect 293092 335656 293098 335668
rect 293678 335656 293684 335668
rect 293736 335656 293742 335708
rect 296806 335656 296812 335708
rect 296864 335696 296870 335708
rect 297450 335696 297456 335708
rect 296864 335668 297456 335696
rect 296864 335656 296870 335668
rect 297450 335656 297456 335668
rect 297508 335656 297514 335708
rect 307754 335656 307760 335708
rect 307812 335696 307818 335708
rect 308582 335696 308588 335708
rect 307812 335668 308588 335696
rect 307812 335656 307818 335668
rect 308582 335656 308588 335668
rect 308640 335656 308646 335708
rect 310974 335656 310980 335708
rect 311032 335696 311038 335708
rect 311710 335696 311716 335708
rect 311032 335668 311716 335696
rect 311032 335656 311038 335668
rect 311710 335656 311716 335668
rect 311768 335656 311774 335708
rect 313642 335656 313648 335708
rect 313700 335696 313706 335708
rect 314194 335696 314200 335708
rect 313700 335668 314200 335696
rect 313700 335656 313706 335668
rect 314194 335656 314200 335668
rect 314252 335656 314258 335708
rect 314746 335656 314752 335708
rect 314804 335696 314810 335708
rect 315850 335696 315856 335708
rect 314804 335668 315856 335696
rect 314804 335656 314810 335668
rect 315850 335656 315856 335668
rect 315908 335656 315914 335708
rect 324314 335656 324320 335708
rect 324372 335696 324378 335708
rect 325050 335696 325056 335708
rect 324372 335668 325056 335696
rect 324372 335656 324378 335668
rect 325050 335656 325056 335668
rect 325108 335656 325114 335708
rect 325786 335656 325792 335708
rect 325844 335696 325850 335708
rect 326246 335696 326252 335708
rect 325844 335668 326252 335696
rect 325844 335656 325850 335668
rect 326246 335656 326252 335668
rect 326304 335656 326310 335708
rect 328454 335656 328460 335708
rect 328512 335696 328518 335708
rect 329006 335696 329012 335708
rect 328512 335668 329012 335696
rect 328512 335656 328518 335668
rect 329006 335656 329012 335668
rect 329064 335656 329070 335708
rect 338298 335656 338304 335708
rect 338356 335696 338362 335708
rect 338758 335696 338764 335708
rect 338356 335668 338764 335696
rect 338356 335656 338362 335668
rect 338758 335656 338764 335668
rect 338816 335656 338822 335708
rect 339494 335656 339500 335708
rect 339552 335696 339558 335708
rect 339954 335696 339960 335708
rect 339552 335668 339960 335696
rect 339552 335656 339558 335668
rect 339954 335656 339960 335668
rect 340012 335656 340018 335708
rect 342714 335656 342720 335708
rect 342772 335696 342778 335708
rect 342898 335696 342904 335708
rect 342772 335668 342904 335696
rect 342772 335656 342778 335668
rect 342898 335656 342904 335668
rect 342956 335656 342962 335708
rect 345198 335656 345204 335708
rect 345256 335696 345262 335708
rect 346118 335696 346124 335708
rect 345256 335668 346124 335696
rect 345256 335656 345262 335668
rect 346118 335656 346124 335668
rect 346176 335656 346182 335708
rect 348050 335656 348056 335708
rect 348108 335696 348114 335708
rect 348326 335696 348332 335708
rect 348108 335668 348332 335696
rect 348108 335656 348114 335668
rect 348326 335656 348332 335668
rect 348384 335656 348390 335708
rect 229186 335588 229192 335640
rect 229244 335628 229250 335640
rect 230106 335628 230112 335640
rect 229244 335600 230112 335628
rect 229244 335588 229250 335600
rect 230106 335588 230112 335600
rect 230164 335588 230170 335640
rect 231946 335588 231952 335640
rect 232004 335628 232010 335640
rect 232222 335628 232228 335640
rect 232004 335600 232228 335628
rect 232004 335588 232010 335600
rect 232222 335588 232228 335600
rect 232280 335588 232286 335640
rect 233234 335588 233240 335640
rect 233292 335628 233298 335640
rect 233510 335628 233516 335640
rect 233292 335600 233516 335628
rect 233292 335588 233298 335600
rect 233510 335588 233516 335600
rect 233568 335588 233574 335640
rect 234706 335588 234712 335640
rect 234764 335628 234770 335640
rect 234982 335628 234988 335640
rect 234764 335600 234988 335628
rect 234764 335588 234770 335600
rect 234982 335588 234988 335600
rect 235040 335588 235046 335640
rect 235166 335588 235172 335640
rect 235224 335628 235230 335640
rect 235718 335628 235724 335640
rect 235224 335600 235724 335628
rect 235224 335588 235230 335600
rect 235718 335588 235724 335600
rect 235776 335588 235782 335640
rect 237466 335588 237472 335640
rect 237524 335628 237530 335640
rect 237926 335628 237932 335640
rect 237524 335600 237932 335628
rect 237524 335588 237530 335600
rect 237926 335588 237932 335600
rect 237984 335588 237990 335640
rect 239122 335588 239128 335640
rect 239180 335628 239186 335640
rect 239858 335628 239864 335640
rect 239180 335600 239864 335628
rect 239180 335588 239186 335600
rect 239858 335588 239864 335600
rect 239916 335588 239922 335640
rect 240410 335588 240416 335640
rect 240468 335628 240474 335640
rect 241054 335628 241060 335640
rect 240468 335600 241060 335628
rect 240468 335588 240474 335600
rect 241054 335588 241060 335600
rect 241112 335588 241118 335640
rect 241606 335588 241612 335640
rect 241664 335628 241670 335640
rect 242342 335628 242348 335640
rect 241664 335600 242348 335628
rect 241664 335588 241670 335600
rect 242342 335588 242348 335600
rect 242400 335588 242406 335640
rect 244274 335588 244280 335640
rect 244332 335628 244338 335640
rect 245194 335628 245200 335640
rect 244332 335600 245200 335628
rect 244332 335588 244338 335600
rect 245194 335588 245200 335600
rect 245252 335588 245258 335640
rect 247494 335588 247500 335640
rect 247552 335628 247558 335640
rect 247954 335628 247960 335640
rect 247552 335600 247960 335628
rect 247552 335588 247558 335600
rect 247954 335588 247960 335600
rect 248012 335588 248018 335640
rect 248690 335588 248696 335640
rect 248748 335628 248754 335640
rect 249426 335628 249432 335640
rect 248748 335600 249432 335628
rect 248748 335588 248754 335600
rect 249426 335588 249432 335600
rect 249484 335588 249490 335640
rect 250162 335588 250168 335640
rect 250220 335628 250226 335640
rect 250898 335628 250904 335640
rect 250220 335600 250904 335628
rect 250220 335588 250226 335600
rect 250898 335588 250904 335600
rect 250956 335588 250962 335640
rect 251634 335588 251640 335640
rect 251692 335628 251698 335640
rect 252094 335628 252100 335640
rect 251692 335600 252100 335628
rect 251692 335588 251698 335600
rect 252094 335588 252100 335600
rect 252152 335588 252158 335640
rect 252554 335588 252560 335640
rect 252612 335628 252618 335640
rect 253106 335628 253112 335640
rect 252612 335600 253112 335628
rect 252612 335588 252618 335600
rect 253106 335588 253112 335600
rect 253164 335588 253170 335640
rect 254118 335588 254124 335640
rect 254176 335628 254182 335640
rect 254762 335628 254768 335640
rect 254176 335600 254768 335628
rect 254176 335588 254182 335600
rect 254762 335588 254768 335600
rect 254820 335588 254826 335640
rect 255774 335588 255780 335640
rect 255832 335628 255838 335640
rect 256234 335628 256240 335640
rect 255832 335600 256240 335628
rect 255832 335588 255838 335600
rect 256234 335588 256240 335600
rect 256292 335588 256298 335640
rect 257338 335588 257344 335640
rect 257396 335628 257402 335640
rect 257706 335628 257712 335640
rect 257396 335600 257712 335628
rect 257396 335588 257402 335600
rect 257706 335588 257712 335600
rect 257764 335588 257770 335640
rect 258626 335588 258632 335640
rect 258684 335628 258690 335640
rect 259178 335628 259184 335640
rect 258684 335600 259184 335628
rect 258684 335588 258690 335600
rect 259178 335588 259184 335600
rect 259236 335588 259242 335640
rect 259638 335588 259644 335640
rect 259696 335628 259702 335640
rect 260374 335628 260380 335640
rect 259696 335600 260380 335628
rect 259696 335588 259702 335600
rect 260374 335588 260380 335600
rect 260432 335588 260438 335640
rect 261202 335588 261208 335640
rect 261260 335628 261266 335640
rect 261662 335628 261668 335640
rect 261260 335600 261668 335628
rect 261260 335588 261266 335600
rect 261662 335588 261668 335600
rect 261720 335588 261726 335640
rect 262398 335588 262404 335640
rect 262456 335628 262462 335640
rect 262674 335628 262680 335640
rect 262456 335600 262680 335628
rect 262456 335588 262462 335600
rect 262674 335588 262680 335600
rect 262732 335588 262738 335640
rect 263962 335588 263968 335640
rect 264020 335628 264026 335640
rect 264882 335628 264888 335640
rect 264020 335600 264888 335628
rect 264020 335588 264026 335600
rect 264882 335588 264888 335600
rect 264940 335588 264946 335640
rect 265158 335588 265164 335640
rect 265216 335628 265222 335640
rect 265342 335628 265348 335640
rect 265216 335600 265348 335628
rect 265216 335588 265222 335600
rect 265342 335588 265348 335600
rect 265400 335588 265406 335640
rect 266354 335588 266360 335640
rect 266412 335628 266418 335640
rect 266814 335628 266820 335640
rect 266412 335600 266820 335628
rect 266412 335588 266418 335600
rect 266814 335588 266820 335600
rect 266872 335588 266878 335640
rect 268378 335588 268384 335640
rect 268436 335628 268442 335640
rect 269022 335628 269028 335640
rect 268436 335600 269028 335628
rect 268436 335588 268442 335600
rect 269022 335588 269028 335600
rect 269080 335588 269086 335640
rect 269666 335588 269672 335640
rect 269724 335628 269730 335640
rect 270402 335628 270408 335640
rect 269724 335600 270408 335628
rect 269724 335588 269730 335600
rect 270402 335588 270408 335600
rect 270460 335588 270466 335640
rect 270494 335588 270500 335640
rect 270552 335628 270558 335640
rect 271598 335628 271604 335640
rect 270552 335600 271604 335628
rect 270552 335588 270558 335600
rect 271598 335588 271604 335600
rect 271656 335588 271662 335640
rect 272058 335588 272064 335640
rect 272116 335628 272122 335640
rect 273162 335628 273168 335640
rect 272116 335600 273168 335628
rect 272116 335588 272122 335600
rect 273162 335588 273168 335600
rect 273220 335588 273226 335640
rect 273714 335588 273720 335640
rect 273772 335628 273778 335640
rect 274542 335628 274548 335640
rect 273772 335600 274548 335628
rect 273772 335588 273778 335600
rect 274542 335588 274548 335600
rect 274600 335588 274606 335640
rect 276106 335588 276112 335640
rect 276164 335628 276170 335640
rect 276566 335628 276572 335640
rect 276164 335600 276572 335628
rect 276164 335588 276170 335600
rect 276566 335588 276572 335600
rect 276624 335588 276630 335640
rect 277762 335588 277768 335640
rect 277820 335628 277826 335640
rect 278314 335628 278320 335640
rect 277820 335600 278320 335628
rect 277820 335588 277826 335600
rect 278314 335588 278320 335600
rect 278372 335588 278378 335640
rect 280338 335588 280344 335640
rect 280396 335628 280402 335640
rect 280706 335628 280712 335640
rect 280396 335600 280712 335628
rect 280396 335588 280402 335600
rect 280706 335588 280712 335600
rect 280764 335588 280770 335640
rect 282270 335588 282276 335640
rect 282328 335628 282334 335640
rect 282822 335628 282828 335640
rect 282328 335600 282828 335628
rect 282328 335588 282334 335600
rect 282822 335588 282828 335600
rect 282880 335588 282886 335640
rect 283282 335588 283288 335640
rect 283340 335628 283346 335640
rect 283926 335628 283932 335640
rect 283340 335600 283932 335628
rect 283340 335588 283346 335600
rect 283926 335588 283932 335600
rect 283984 335588 283990 335640
rect 285674 335588 285680 335640
rect 285732 335628 285738 335640
rect 286410 335628 286416 335640
rect 285732 335600 286416 335628
rect 285732 335588 285738 335600
rect 286410 335588 286416 335600
rect 286468 335588 286474 335640
rect 287606 335588 287612 335640
rect 287664 335628 287670 335640
rect 288066 335628 288072 335640
rect 287664 335600 288072 335628
rect 287664 335588 287670 335600
rect 288066 335588 288072 335600
rect 288124 335588 288130 335640
rect 288526 335588 288532 335640
rect 288584 335628 288590 335640
rect 289078 335628 289084 335640
rect 288584 335600 289084 335628
rect 288584 335588 288590 335600
rect 289078 335588 289084 335600
rect 289136 335588 289142 335640
rect 289814 335588 289820 335640
rect 289872 335628 289878 335640
rect 290550 335628 290556 335640
rect 289872 335600 290556 335628
rect 289872 335588 289878 335600
rect 290550 335588 290556 335600
rect 290608 335588 290614 335640
rect 291470 335588 291476 335640
rect 291528 335628 291534 335640
rect 291838 335628 291844 335640
rect 291528 335600 291844 335628
rect 291528 335588 291534 335600
rect 291838 335588 291844 335600
rect 291896 335588 291902 335640
rect 292942 335588 292948 335640
rect 293000 335628 293006 335640
rect 293494 335628 293500 335640
rect 293000 335600 293500 335628
rect 293000 335588 293006 335600
rect 293494 335588 293500 335600
rect 293552 335588 293558 335640
rect 298462 335588 298468 335640
rect 298520 335628 298526 335640
rect 299106 335628 299112 335640
rect 298520 335600 299112 335628
rect 298520 335588 298526 335600
rect 299106 335588 299112 335600
rect 299164 335588 299170 335640
rect 302602 335588 302608 335640
rect 302660 335628 302666 335640
rect 303430 335628 303436 335640
rect 302660 335600 303436 335628
rect 302660 335588 302666 335600
rect 303430 335588 303436 335600
rect 303488 335588 303494 335640
rect 303982 335588 303988 335640
rect 304040 335628 304046 335640
rect 304534 335628 304540 335640
rect 304040 335600 304540 335628
rect 304040 335588 304046 335600
rect 304534 335588 304540 335600
rect 304592 335588 304598 335640
rect 305178 335588 305184 335640
rect 305236 335628 305242 335640
rect 305730 335628 305736 335640
rect 305236 335600 305736 335628
rect 305236 335588 305242 335600
rect 305730 335588 305736 335600
rect 305788 335588 305794 335640
rect 306650 335588 306656 335640
rect 306708 335628 306714 335640
rect 306926 335628 306932 335640
rect 306708 335600 306932 335628
rect 306708 335588 306714 335600
rect 306926 335588 306932 335600
rect 306984 335588 306990 335640
rect 307938 335588 307944 335640
rect 307996 335628 308002 335640
rect 308674 335628 308680 335640
rect 307996 335600 308680 335628
rect 307996 335588 308002 335600
rect 308674 335588 308680 335600
rect 308732 335588 308738 335640
rect 310514 335588 310520 335640
rect 310572 335628 310578 335640
rect 310698 335628 310704 335640
rect 310572 335600 310704 335628
rect 310572 335588 310578 335600
rect 310698 335588 310704 335600
rect 310756 335588 310762 335640
rect 312170 335588 312176 335640
rect 312228 335628 312234 335640
rect 313182 335628 313188 335640
rect 312228 335600 313188 335628
rect 312228 335588 312234 335600
rect 313182 335588 313188 335600
rect 313240 335588 313246 335640
rect 313274 335588 313280 335640
rect 313332 335628 313338 335640
rect 314286 335628 314292 335640
rect 313332 335600 314292 335628
rect 313332 335588 313338 335600
rect 314286 335588 314292 335600
rect 314344 335588 314350 335640
rect 316126 335588 316132 335640
rect 316184 335628 316190 335640
rect 316954 335628 316960 335640
rect 316184 335600 316960 335628
rect 316184 335588 316190 335600
rect 316954 335588 316960 335600
rect 317012 335588 317018 335640
rect 318978 335588 318984 335640
rect 319036 335628 319042 335640
rect 319438 335628 319444 335640
rect 319036 335600 319444 335628
rect 319036 335588 319042 335600
rect 319438 335588 319444 335600
rect 319496 335588 319502 335640
rect 320634 335588 320640 335640
rect 320692 335628 320698 335640
rect 321094 335628 321100 335640
rect 320692 335600 321100 335628
rect 320692 335588 320698 335600
rect 321094 335588 321100 335600
rect 321152 335588 321158 335640
rect 324774 335588 324780 335640
rect 324832 335628 324838 335640
rect 325326 335628 325332 335640
rect 324832 335600 325332 335628
rect 324832 335588 324838 335600
rect 325326 335588 325332 335600
rect 325384 335588 325390 335640
rect 325878 335588 325884 335640
rect 325936 335628 325942 335640
rect 326338 335628 326344 335640
rect 325936 335600 326344 335628
rect 325936 335588 325942 335600
rect 326338 335588 326344 335600
rect 326396 335588 326402 335640
rect 327258 335588 327264 335640
rect 327316 335628 327322 335640
rect 327534 335628 327540 335640
rect 327316 335600 327540 335628
rect 327316 335588 327322 335600
rect 327534 335588 327540 335600
rect 327592 335588 327598 335640
rect 329926 335588 329932 335640
rect 329984 335628 329990 335640
rect 330478 335628 330484 335640
rect 329984 335600 330484 335628
rect 329984 335588 329990 335600
rect 330478 335588 330484 335600
rect 330536 335588 330542 335640
rect 331398 335588 331404 335640
rect 331456 335628 331462 335640
rect 332134 335628 332140 335640
rect 331456 335600 332140 335628
rect 331456 335588 331462 335600
rect 332134 335588 332140 335600
rect 332192 335588 332198 335640
rect 332686 335588 332692 335640
rect 332744 335628 332750 335640
rect 333422 335628 333428 335640
rect 332744 335600 333428 335628
rect 332744 335588 332750 335600
rect 333422 335588 333428 335600
rect 333480 335588 333486 335640
rect 334342 335588 334348 335640
rect 334400 335628 334406 335640
rect 334618 335628 334624 335640
rect 334400 335600 334624 335628
rect 334400 335588 334406 335600
rect 334618 335588 334624 335600
rect 334676 335588 334682 335640
rect 337010 335588 337016 335640
rect 337068 335628 337074 335640
rect 337562 335628 337568 335640
rect 337068 335600 337568 335628
rect 337068 335588 337074 335600
rect 337562 335588 337568 335600
rect 337620 335588 337626 335640
rect 338482 335588 338488 335640
rect 338540 335628 338546 335640
rect 339034 335628 339040 335640
rect 338540 335600 339040 335628
rect 338540 335588 338546 335600
rect 339034 335588 339040 335600
rect 339092 335588 339098 335640
rect 339770 335588 339776 335640
rect 339828 335628 339834 335640
rect 340506 335628 340512 335640
rect 339828 335600 340512 335628
rect 339828 335588 339834 335600
rect 340506 335588 340512 335600
rect 340564 335588 340570 335640
rect 340966 335588 340972 335640
rect 341024 335628 341030 335640
rect 341702 335628 341708 335640
rect 341024 335600 341708 335628
rect 341024 335588 341030 335600
rect 341702 335588 341708 335600
rect 341760 335588 341766 335640
rect 342438 335588 342444 335640
rect 342496 335628 342502 335640
rect 343174 335628 343180 335640
rect 342496 335600 343180 335628
rect 342496 335588 342502 335600
rect 343174 335588 343180 335600
rect 343232 335588 343238 335640
rect 343910 335588 343916 335640
rect 343968 335628 343974 335640
rect 344186 335628 344192 335640
rect 343968 335600 344192 335628
rect 343968 335588 343974 335600
rect 344186 335588 344192 335600
rect 344244 335588 344250 335640
rect 345014 335588 345020 335640
rect 345072 335628 345078 335640
rect 345658 335628 345664 335640
rect 345072 335600 345664 335628
rect 345072 335588 345078 335600
rect 345658 335588 345664 335600
rect 345716 335588 345722 335640
rect 347774 335588 347780 335640
rect 347832 335628 347838 335640
rect 348418 335628 348424 335640
rect 347832 335600 348424 335628
rect 347832 335588 347838 335600
rect 348418 335588 348424 335600
rect 348476 335588 348482 335640
rect 248506 335520 248512 335572
rect 248564 335560 248570 335572
rect 249150 335560 249156 335572
rect 248564 335532 249156 335560
rect 248564 335520 248570 335532
rect 249150 335520 249156 335532
rect 249208 335520 249214 335572
rect 249978 335520 249984 335572
rect 250036 335560 250042 335572
rect 250622 335560 250628 335572
rect 250036 335532 250628 335560
rect 250036 335520 250042 335532
rect 250622 335520 250628 335532
rect 250680 335520 250686 335572
rect 251450 335520 251456 335572
rect 251508 335560 251514 335572
rect 252370 335560 252376 335572
rect 251508 335532 252376 335560
rect 251508 335520 251514 335532
rect 252370 335520 252376 335532
rect 252428 335520 252434 335572
rect 277578 335520 277584 335572
rect 277636 335560 277642 335572
rect 278498 335560 278504 335572
rect 277636 335532 278504 335560
rect 277636 335520 277642 335532
rect 278498 335520 278504 335532
rect 278556 335520 278562 335572
rect 287146 335520 287152 335572
rect 287204 335560 287210 335572
rect 287974 335560 287980 335572
rect 287204 335532 287980 335560
rect 287204 335520 287210 335532
rect 287974 335520 287980 335532
rect 288032 335520 288038 335572
rect 291286 335520 291292 335572
rect 291344 335560 291350 335572
rect 292206 335560 292212 335572
rect 291344 335532 292212 335560
rect 291344 335520 291350 335532
rect 292206 335520 292212 335532
rect 292264 335520 292270 335572
rect 292758 335520 292764 335572
rect 292816 335560 292822 335572
rect 293402 335560 293408 335572
rect 292816 335532 293408 335560
rect 292816 335520 292822 335532
rect 293402 335520 293408 335532
rect 293460 335520 293466 335572
rect 312078 335520 312084 335572
rect 312136 335560 312142 335572
rect 312630 335560 312636 335572
rect 312136 335532 312636 335560
rect 312136 335520 312142 335532
rect 312630 335520 312636 335532
rect 312688 335520 312694 335572
rect 317782 335520 317788 335572
rect 317840 335560 317846 335572
rect 318058 335560 318064 335572
rect 317840 335532 318064 335560
rect 317840 335520 317846 335532
rect 318058 335520 318064 335532
rect 318116 335520 318122 335572
rect 345106 335520 345112 335572
rect 345164 335560 345170 335572
rect 345382 335560 345388 335572
rect 345164 335532 345388 335560
rect 345164 335520 345170 335532
rect 345382 335520 345388 335532
rect 345440 335520 345446 335572
rect 233510 335452 233516 335504
rect 233568 335492 233574 335504
rect 233970 335492 233976 335504
rect 233568 335464 233976 335492
rect 233568 335452 233574 335464
rect 233970 335452 233976 335464
rect 234028 335452 234034 335504
rect 234982 335452 234988 335504
rect 235040 335492 235046 335504
rect 235442 335492 235448 335504
rect 235040 335464 235448 335492
rect 235040 335452 235046 335464
rect 235442 335452 235448 335464
rect 235500 335452 235506 335504
rect 243078 335452 243084 335504
rect 243136 335492 243142 335504
rect 243998 335492 244004 335504
rect 243136 335464 244004 335492
rect 243136 335452 243142 335464
rect 243998 335452 244004 335464
rect 244056 335452 244062 335504
rect 258166 335452 258172 335504
rect 258224 335492 258230 335504
rect 258994 335492 259000 335504
rect 258224 335464 259000 335492
rect 258224 335452 258230 335464
rect 258994 335452 259000 335464
rect 259052 335452 259058 335504
rect 262398 335452 262404 335504
rect 262456 335492 262462 335504
rect 263134 335492 263140 335504
rect 262456 335464 263140 335492
rect 262456 335452 262462 335464
rect 263134 335452 263140 335464
rect 263192 335452 263198 335504
rect 266814 335452 266820 335504
rect 266872 335492 266878 335504
rect 267366 335492 267372 335504
rect 266872 335464 267372 335492
rect 266872 335452 266878 335464
rect 267366 335452 267372 335464
rect 267424 335452 267430 335504
rect 276106 335452 276112 335504
rect 276164 335492 276170 335504
rect 276658 335492 276664 335504
rect 276164 335464 276664 335492
rect 276164 335452 276170 335464
rect 276658 335452 276664 335464
rect 276716 335452 276722 335504
rect 311066 335452 311072 335504
rect 311124 335492 311130 335504
rect 311618 335492 311624 335504
rect 311124 335464 311624 335492
rect 311124 335452 311130 335464
rect 311618 335452 311624 335464
rect 311676 335452 311682 335504
rect 315022 335452 315028 335504
rect 315080 335492 315086 335504
rect 315298 335492 315304 335504
rect 315080 335464 315304 335492
rect 315080 335452 315086 335464
rect 315298 335452 315304 335464
rect 315356 335452 315362 335504
rect 327350 335452 327356 335504
rect 327408 335492 327414 335504
rect 327534 335492 327540 335504
rect 327408 335464 327540 335492
rect 327408 335452 327414 335464
rect 327534 335452 327540 335464
rect 327592 335452 327598 335504
rect 342530 335452 342536 335504
rect 342588 335492 342594 335504
rect 343450 335492 343456 335504
rect 342588 335464 343456 335492
rect 342588 335452 342594 335464
rect 343450 335452 343456 335464
rect 343508 335452 343514 335504
rect 238846 335384 238852 335436
rect 238904 335424 238910 335436
rect 239214 335424 239220 335436
rect 238904 335396 239220 335424
rect 238904 335384 238910 335396
rect 239214 335384 239220 335396
rect 239272 335384 239278 335436
rect 258626 335384 258632 335436
rect 258684 335424 258690 335436
rect 259270 335424 259276 335436
rect 258684 335396 259276 335424
rect 258684 335384 258690 335396
rect 259270 335384 259276 335396
rect 259328 335384 259334 335436
rect 320910 335384 320916 335436
rect 320968 335424 320974 335436
rect 321462 335424 321468 335436
rect 320968 335396 321468 335424
rect 320968 335384 320974 335396
rect 321462 335384 321468 335396
rect 321520 335384 321526 335436
rect 296990 335316 296996 335368
rect 297048 335356 297054 335368
rect 297910 335356 297916 335368
rect 297048 335328 297916 335356
rect 297048 335316 297054 335328
rect 297910 335316 297916 335328
rect 297968 335316 297974 335368
rect 327350 335316 327356 335368
rect 327408 335356 327414 335368
rect 328270 335356 328276 335368
rect 327408 335328 328276 335356
rect 327408 335316 327414 335328
rect 328270 335316 328276 335328
rect 328328 335316 328334 335368
rect 238846 335248 238852 335300
rect 238904 335288 238910 335300
rect 239582 335288 239588 335300
rect 238904 335260 239588 335288
rect 238904 335248 238910 335260
rect 239582 335248 239588 335260
rect 239640 335248 239646 335300
rect 269758 335180 269764 335232
rect 269816 335220 269822 335232
rect 270126 335220 270132 335232
rect 269816 335192 270132 335220
rect 269816 335180 269822 335192
rect 270126 335180 270132 335192
rect 270184 335180 270190 335232
rect 320174 335180 320180 335232
rect 320232 335220 320238 335232
rect 320269 335223 320327 335229
rect 320269 335220 320281 335223
rect 320232 335192 320281 335220
rect 320232 335180 320238 335192
rect 320269 335189 320281 335192
rect 320315 335189 320327 335223
rect 320269 335183 320327 335189
rect 325878 335180 325884 335232
rect 325936 335220 325942 335232
rect 326522 335220 326528 335232
rect 325936 335192 326528 335220
rect 325936 335180 325942 335192
rect 326522 335180 326528 335192
rect 326580 335180 326586 335232
rect 265066 334976 265072 335028
rect 265124 335016 265130 335028
rect 266170 335016 266176 335028
rect 265124 334988 266176 335016
rect 265124 334976 265130 334988
rect 266170 334976 266176 334988
rect 266228 334976 266234 335028
rect 323302 334976 323308 335028
rect 323360 335016 323366 335028
rect 324038 335016 324044 335028
rect 323360 334988 324044 335016
rect 323360 334976 323366 334988
rect 324038 334976 324044 334988
rect 324096 334976 324102 335028
rect 275646 334704 275652 334756
rect 275704 334744 275710 334756
rect 275830 334744 275836 334756
rect 275704 334716 275836 334744
rect 275704 334704 275710 334716
rect 275830 334704 275836 334716
rect 275888 334704 275894 334756
rect 278774 334704 278780 334756
rect 278832 334744 278838 334756
rect 279234 334744 279240 334756
rect 278832 334716 279240 334744
rect 278832 334704 278838 334716
rect 279234 334704 279240 334716
rect 279292 334704 279298 334756
rect 333054 334636 333060 334688
rect 333112 334676 333118 334688
rect 333238 334676 333244 334688
rect 333112 334648 333244 334676
rect 333112 334636 333118 334648
rect 333238 334636 333244 334648
rect 333296 334636 333302 334688
rect 244461 334475 244519 334481
rect 244461 334441 244473 334475
rect 244507 334472 244519 334475
rect 244550 334472 244556 334484
rect 244507 334444 244556 334472
rect 244507 334441 244519 334444
rect 244461 334435 244519 334441
rect 244550 334432 244556 334444
rect 244608 334432 244614 334484
rect 256694 334092 256700 334144
rect 256752 334132 256758 334144
rect 257246 334132 257252 334144
rect 256752 334104 257252 334132
rect 256752 334092 256758 334104
rect 257246 334092 257252 334104
rect 257304 334092 257310 334144
rect 336826 333888 336832 333940
rect 336884 333928 336890 333940
rect 337286 333928 337292 333940
rect 336884 333900 337292 333928
rect 336884 333888 336890 333900
rect 337286 333888 337292 333900
rect 337344 333888 337350 333940
rect 336826 333752 336832 333804
rect 336884 333792 336890 333804
rect 337378 333792 337384 333804
rect 336884 333764 337384 333792
rect 336884 333752 336890 333764
rect 337378 333752 337384 333764
rect 337436 333752 337442 333804
rect 262766 333724 262772 333736
rect 262727 333696 262772 333724
rect 262766 333684 262772 333696
rect 262824 333684 262830 333736
rect 288618 333548 288624 333600
rect 288676 333588 288682 333600
rect 289170 333588 289176 333600
rect 288676 333560 289176 333588
rect 288676 333548 288682 333560
rect 289170 333548 289176 333560
rect 289228 333548 289234 333600
rect 274910 333480 274916 333532
rect 274968 333520 274974 333532
rect 275186 333520 275192 333532
rect 274968 333492 275192 333520
rect 274968 333480 274974 333492
rect 275186 333480 275192 333492
rect 275244 333480 275250 333532
rect 288894 333480 288900 333532
rect 288952 333520 288958 333532
rect 289538 333520 289544 333532
rect 288952 333492 289544 333520
rect 288952 333480 288958 333492
rect 289538 333480 289544 333492
rect 289596 333480 289602 333532
rect 261110 333276 261116 333328
rect 261168 333316 261174 333328
rect 261386 333316 261392 333328
rect 261168 333288 261392 333316
rect 261168 333276 261174 333288
rect 261386 333276 261392 333288
rect 261444 333276 261450 333328
rect 293954 333276 293960 333328
rect 294012 333316 294018 333328
rect 295058 333316 295064 333328
rect 294012 333288 295064 333316
rect 294012 333276 294018 333288
rect 295058 333276 295064 333288
rect 295116 333276 295122 333328
rect 306742 333276 306748 333328
rect 306800 333316 306806 333328
rect 307478 333316 307484 333328
rect 306800 333288 307484 333316
rect 306800 333276 306806 333288
rect 307478 333276 307484 333288
rect 307536 333276 307542 333328
rect 261386 333140 261392 333192
rect 261444 333180 261450 333192
rect 261846 333180 261852 333192
rect 261444 333152 261852 333180
rect 261444 333140 261450 333152
rect 261846 333140 261852 333152
rect 261904 333140 261910 333192
rect 294230 333140 294236 333192
rect 294288 333180 294294 333192
rect 294414 333180 294420 333192
rect 294288 333152 294420 333180
rect 294288 333140 294294 333152
rect 294414 333140 294420 333152
rect 294472 333140 294478 333192
rect 308122 332936 308128 332988
rect 308180 332976 308186 332988
rect 308858 332976 308864 332988
rect 308180 332948 308864 332976
rect 308180 332936 308186 332948
rect 308858 332936 308864 332948
rect 308916 332936 308922 332988
rect 298094 332732 298100 332784
rect 298152 332772 298158 332784
rect 298738 332772 298744 332784
rect 298152 332744 298744 332772
rect 298152 332732 298158 332744
rect 298738 332732 298744 332744
rect 298796 332732 298802 332784
rect 236730 332664 236736 332716
rect 236788 332704 236794 332716
rect 237190 332704 237196 332716
rect 236788 332676 237196 332704
rect 236788 332664 236794 332676
rect 237190 332664 237196 332676
rect 237248 332664 237254 332716
rect 283006 332664 283012 332716
rect 283064 332704 283070 332716
rect 283466 332704 283472 332716
rect 283064 332676 283472 332704
rect 283064 332664 283070 332676
rect 283466 332664 283472 332676
rect 283524 332664 283530 332716
rect 263870 332324 263876 332376
rect 263928 332364 263934 332376
rect 264698 332364 264704 332376
rect 263928 332336 264704 332364
rect 263928 332324 263934 332336
rect 264698 332324 264704 332336
rect 264756 332324 264762 332376
rect 326062 332256 326068 332308
rect 326120 332296 326126 332308
rect 326798 332296 326804 332308
rect 326120 332268 326804 332296
rect 326120 332256 326126 332268
rect 326798 332256 326804 332268
rect 326856 332256 326862 332308
rect 246206 332052 246212 332104
rect 246264 332092 246270 332104
rect 246666 332092 246672 332104
rect 246264 332064 246672 332092
rect 246264 332052 246270 332064
rect 246666 332052 246672 332064
rect 246724 332052 246730 332104
rect 287330 332052 287336 332104
rect 287388 332092 287394 332104
rect 287882 332092 287888 332104
rect 287388 332064 287888 332092
rect 287388 332052 287394 332064
rect 287882 332052 287888 332064
rect 287940 332052 287946 332104
rect 241882 331984 241888 332036
rect 241940 332024 241946 332036
rect 242158 332024 242164 332036
rect 241940 331996 242164 332024
rect 241940 331984 241946 331996
rect 242158 331984 242164 331996
rect 242216 331984 242222 332036
rect 231026 331848 231032 331900
rect 231084 331888 231090 331900
rect 231302 331888 231308 331900
rect 231084 331860 231308 331888
rect 231084 331848 231090 331860
rect 231302 331848 231308 331860
rect 231360 331848 231366 331900
rect 272242 331848 272248 331900
rect 272300 331888 272306 331900
rect 273070 331888 273076 331900
rect 272300 331860 273076 331888
rect 272300 331848 272306 331860
rect 273070 331848 273076 331860
rect 273128 331848 273134 331900
rect 311250 331848 311256 331900
rect 311308 331888 311314 331900
rect 311434 331888 311440 331900
rect 311308 331860 311440 331888
rect 311308 331848 311314 331860
rect 311434 331848 311440 331860
rect 311492 331848 311498 331900
rect 329006 331848 329012 331900
rect 329064 331888 329070 331900
rect 329558 331888 329564 331900
rect 329064 331860 329564 331888
rect 329064 331848 329070 331860
rect 329558 331848 329564 331860
rect 329616 331848 329622 331900
rect 333238 331848 333244 331900
rect 333296 331888 333302 331900
rect 333698 331888 333704 331900
rect 333296 331860 333704 331888
rect 333296 331848 333302 331860
rect 333698 331848 333704 331860
rect 333756 331848 333762 331900
rect 323394 331712 323400 331764
rect 323452 331752 323458 331764
rect 323854 331752 323860 331764
rect 323452 331724 323860 331752
rect 323452 331712 323458 331724
rect 323854 331712 323860 331724
rect 323912 331712 323918 331764
rect 298186 331372 298192 331424
rect 298244 331412 298250 331424
rect 298830 331412 298836 331424
rect 298244 331384 298836 331412
rect 298244 331372 298250 331384
rect 298830 331372 298836 331384
rect 298888 331372 298894 331424
rect 301222 331304 301228 331356
rect 301280 331304 301286 331356
rect 240778 331276 240784 331288
rect 240704 331248 240784 331276
rect 240704 331016 240732 331248
rect 240778 331236 240784 331248
rect 240836 331236 240842 331288
rect 245838 331236 245844 331288
rect 245896 331236 245902 331288
rect 260190 331276 260196 331288
rect 260024 331248 260196 331276
rect 245856 331140 245884 331236
rect 260024 331220 260052 331248
rect 260190 331236 260196 331248
rect 260248 331236 260254 331288
rect 260006 331168 260012 331220
rect 260064 331168 260070 331220
rect 246022 331140 246028 331152
rect 245856 331112 246028 331140
rect 246022 331100 246028 331112
rect 246080 331100 246086 331152
rect 298738 331100 298744 331152
rect 298796 331140 298802 331152
rect 299198 331140 299204 331152
rect 298796 331112 299204 331140
rect 298796 331100 298802 331112
rect 299198 331100 299204 331112
rect 299256 331100 299262 331152
rect 301240 331084 301268 331304
rect 304718 331276 304724 331288
rect 304276 331248 304724 331276
rect 304276 331220 304304 331248
rect 304718 331236 304724 331248
rect 304776 331236 304782 331288
rect 309870 331236 309876 331288
rect 309928 331236 309934 331288
rect 304258 331168 304264 331220
rect 304316 331168 304322 331220
rect 309686 331168 309692 331220
rect 309744 331208 309750 331220
rect 309888 331208 309916 331236
rect 309744 331180 309916 331208
rect 309744 331168 309750 331180
rect 290090 331032 290096 331084
rect 290148 331072 290154 331084
rect 290366 331072 290372 331084
rect 290148 331044 290372 331072
rect 290148 331032 290154 331044
rect 290366 331032 290372 331044
rect 290424 331032 290430 331084
rect 301222 331032 301228 331084
rect 301280 331032 301286 331084
rect 240686 330964 240692 331016
rect 240744 330964 240750 331016
rect 295610 330828 295616 330880
rect 295668 330868 295674 330880
rect 296530 330868 296536 330880
rect 295668 330840 296536 330868
rect 295668 330828 295674 330840
rect 296530 330828 296536 330840
rect 296588 330828 296594 330880
rect 258258 330692 258264 330744
rect 258316 330732 258322 330744
rect 259362 330732 259368 330744
rect 258316 330704 259368 330732
rect 258316 330692 258322 330704
rect 259362 330692 259368 330704
rect 259420 330692 259426 330744
rect 341518 330624 341524 330676
rect 341576 330664 341582 330676
rect 342070 330664 342076 330676
rect 341576 330636 342076 330664
rect 341576 330624 341582 330636
rect 342070 330624 342076 330636
rect 342128 330624 342134 330676
rect 302326 330556 302332 330608
rect 302384 330596 302390 330608
rect 303154 330596 303160 330608
rect 302384 330568 303160 330596
rect 302384 330556 302390 330568
rect 303154 330556 303160 330568
rect 303212 330556 303218 330608
rect 320358 330556 320364 330608
rect 320416 330596 320422 330608
rect 321370 330596 321376 330608
rect 320416 330568 321376 330596
rect 320416 330556 320422 330568
rect 321370 330556 321376 330568
rect 321428 330556 321434 330608
rect 323210 330556 323216 330608
rect 323268 330596 323274 330608
rect 324222 330596 324228 330608
rect 323268 330568 324228 330596
rect 323268 330556 323274 330568
rect 324222 330556 324228 330568
rect 324280 330556 324286 330608
rect 288618 330488 288624 330540
rect 288676 330528 288682 330540
rect 289354 330528 289360 330540
rect 288676 330500 289360 330528
rect 288676 330488 288682 330500
rect 289354 330488 289360 330500
rect 289412 330488 289418 330540
rect 321830 330488 321836 330540
rect 321888 330528 321894 330540
rect 322658 330528 322664 330540
rect 321888 330500 322664 330528
rect 321888 330488 321894 330500
rect 322658 330488 322664 330500
rect 322716 330488 322722 330540
rect 323118 330488 323124 330540
rect 323176 330528 323182 330540
rect 324038 330528 324044 330540
rect 323176 330500 324044 330528
rect 323176 330488 323182 330500
rect 324038 330488 324044 330500
rect 324096 330488 324102 330540
rect 321646 330420 321652 330472
rect 321704 330460 321710 330472
rect 322750 330460 322756 330472
rect 321704 330432 322756 330460
rect 321704 330420 321710 330432
rect 322750 330420 322756 330432
rect 322808 330420 322814 330472
rect 322934 330420 322940 330472
rect 322992 330460 322998 330472
rect 323946 330460 323952 330472
rect 322992 330432 323952 330460
rect 322992 330420 322998 330432
rect 323946 330420 323952 330432
rect 324004 330420 324010 330472
rect 321554 330352 321560 330404
rect 321612 330392 321618 330404
rect 322474 330392 322480 330404
rect 321612 330364 322480 330392
rect 321612 330352 321618 330364
rect 322474 330352 322480 330364
rect 322532 330352 322538 330404
rect 317506 330284 317512 330336
rect 317564 330324 317570 330336
rect 318610 330324 318616 330336
rect 317564 330296 318616 330324
rect 317564 330284 317570 330296
rect 318610 330284 318616 330296
rect 318668 330284 318674 330336
rect 304994 329944 305000 329996
rect 305052 329984 305058 329996
rect 305454 329984 305460 329996
rect 305052 329956 305460 329984
rect 305052 329944 305058 329956
rect 305454 329944 305460 329956
rect 305512 329944 305518 329996
rect 245930 329128 245936 329180
rect 245988 329168 245994 329180
rect 246114 329168 246120 329180
rect 245988 329140 246120 329168
rect 245988 329128 245994 329140
rect 246114 329128 246120 329140
rect 246172 329128 246178 329180
rect 295426 328720 295432 328772
rect 295484 328760 295490 328772
rect 296346 328760 296352 328772
rect 295484 328732 296352 328760
rect 295484 328720 295490 328732
rect 296346 328720 296352 328732
rect 296404 328720 296410 328772
rect 242526 328556 242532 328568
rect 242268 328528 242532 328556
rect 242268 328500 242296 328528
rect 242526 328516 242532 328528
rect 242584 328516 242590 328568
rect 286134 328556 286140 328568
rect 285876 328528 286140 328556
rect 285876 328500 285904 328528
rect 286134 328516 286140 328528
rect 286192 328516 286198 328568
rect 299842 328516 299848 328568
rect 299900 328556 299906 328568
rect 300118 328556 300124 328568
rect 299900 328528 300124 328556
rect 299900 328516 299906 328528
rect 300118 328516 300124 328528
rect 300176 328516 300182 328568
rect 301038 328516 301044 328568
rect 301096 328556 301102 328568
rect 301590 328556 301596 328568
rect 301096 328528 301596 328556
rect 301096 328516 301102 328528
rect 301590 328516 301596 328528
rect 301648 328516 301654 328568
rect 306650 328516 306656 328568
rect 306708 328556 306714 328568
rect 307570 328556 307576 328568
rect 306708 328528 307576 328556
rect 306708 328516 306714 328528
rect 307570 328516 307576 328528
rect 307628 328516 307634 328568
rect 232130 328488 232136 328500
rect 232091 328460 232136 328488
rect 232130 328448 232136 328460
rect 232188 328448 232194 328500
rect 242250 328448 242256 328500
rect 242308 328448 242314 328500
rect 243630 328448 243636 328500
rect 243688 328488 243694 328500
rect 243814 328488 243820 328500
rect 243688 328460 243820 328488
rect 243688 328448 243694 328460
rect 243814 328448 243820 328460
rect 243872 328448 243878 328500
rect 244458 328488 244464 328500
rect 244419 328460 244464 328488
rect 244458 328448 244464 328460
rect 244516 328448 244522 328500
rect 253106 328448 253112 328500
rect 253164 328488 253170 328500
rect 253658 328488 253664 328500
rect 253164 328460 253664 328488
rect 253164 328448 253170 328460
rect 253658 328448 253664 328460
rect 253716 328448 253722 328500
rect 265434 328448 265440 328500
rect 265492 328488 265498 328500
rect 265526 328488 265532 328500
rect 265492 328460 265532 328488
rect 265492 328448 265498 328460
rect 265526 328448 265532 328460
rect 265584 328448 265590 328500
rect 277578 328448 277584 328500
rect 277636 328488 277642 328500
rect 278498 328488 278504 328500
rect 277636 328460 278504 328488
rect 277636 328448 277642 328460
rect 278498 328448 278504 328460
rect 278556 328448 278562 328500
rect 284662 328448 284668 328500
rect 284720 328488 284726 328500
rect 285490 328488 285496 328500
rect 284720 328460 285496 328488
rect 284720 328448 284726 328460
rect 285490 328448 285496 328460
rect 285548 328448 285554 328500
rect 285858 328448 285864 328500
rect 285916 328448 285922 328500
rect 285950 328448 285956 328500
rect 286008 328488 286014 328500
rect 286594 328488 286600 328500
rect 286008 328460 286600 328488
rect 286008 328448 286014 328460
rect 286594 328448 286600 328460
rect 286652 328448 286658 328500
rect 326246 328448 326252 328500
rect 326304 328488 326310 328500
rect 326304 328460 326384 328488
rect 326304 328448 326310 328460
rect 326356 328432 326384 328460
rect 100662 328420 100668 328432
rect 100623 328392 100668 328420
rect 100662 328380 100668 328392
rect 100720 328380 100726 328432
rect 231118 328420 231124 328432
rect 231079 328392 231124 328420
rect 231118 328380 231124 328392
rect 231176 328380 231182 328432
rect 254670 328420 254676 328432
rect 254631 328392 254676 328420
rect 254670 328380 254676 328392
rect 254728 328380 254734 328432
rect 258626 328380 258632 328432
rect 258684 328420 258690 328432
rect 258810 328420 258816 328432
rect 258684 328392 258816 328420
rect 258684 328380 258690 328392
rect 258810 328380 258816 328392
rect 258868 328380 258874 328432
rect 263686 328380 263692 328432
rect 263744 328380 263750 328432
rect 280614 328420 280620 328432
rect 280575 328392 280620 328420
rect 280614 328380 280620 328392
rect 280672 328380 280678 328432
rect 281902 328420 281908 328432
rect 281863 328392 281908 328420
rect 281902 328380 281908 328392
rect 281960 328380 281966 328432
rect 290274 328380 290280 328432
rect 290332 328420 290338 328432
rect 290642 328420 290648 328432
rect 290332 328392 290648 328420
rect 290332 328380 290338 328392
rect 290642 328380 290648 328392
rect 290700 328380 290706 328432
rect 291746 328380 291752 328432
rect 291804 328420 291810 328432
rect 291930 328420 291936 328432
rect 291804 328392 291936 328420
rect 291804 328380 291810 328392
rect 291930 328380 291936 328392
rect 291988 328380 291994 328432
rect 319438 328420 319444 328432
rect 319399 328392 319444 328420
rect 319438 328380 319444 328392
rect 319496 328380 319502 328432
rect 326338 328380 326344 328432
rect 326396 328380 326402 328432
rect 341518 328380 341524 328432
rect 341576 328420 341582 328432
rect 341702 328420 341708 328432
rect 341576 328392 341708 328420
rect 341576 328380 341582 328392
rect 341702 328380 341708 328392
rect 341760 328380 341766 328432
rect 344278 328420 344284 328432
rect 344239 328392 344284 328420
rect 344278 328380 344284 328392
rect 344336 328380 344342 328432
rect 263704 328352 263732 328380
rect 263778 328352 263784 328364
rect 263704 328324 263784 328352
rect 263778 328312 263784 328324
rect 263836 328312 263842 328364
rect 270494 328312 270500 328364
rect 270552 328352 270558 328364
rect 271506 328352 271512 328364
rect 270552 328324 271512 328352
rect 270552 328312 270558 328324
rect 271506 328312 271512 328324
rect 271564 328312 271570 328364
rect 284478 328244 284484 328296
rect 284536 328284 284542 328296
rect 285306 328284 285312 328296
rect 284536 328256 285312 328284
rect 284536 328244 284542 328256
rect 285306 328244 285312 328256
rect 285364 328244 285370 328296
rect 265250 328176 265256 328228
rect 265308 328216 265314 328228
rect 266078 328216 266084 328228
rect 265308 328188 266084 328216
rect 265308 328176 265314 328188
rect 266078 328176 266084 328188
rect 266136 328176 266142 328228
rect 269574 327904 269580 327956
rect 269632 327944 269638 327956
rect 270034 327944 270040 327956
rect 269632 327916 270040 327944
rect 269632 327904 269638 327916
rect 270034 327904 270040 327916
rect 270092 327904 270098 327956
rect 273622 327428 273628 327480
rect 273680 327468 273686 327480
rect 274174 327468 274180 327480
rect 273680 327440 274180 327468
rect 273680 327428 273686 327440
rect 274174 327428 274180 327440
rect 274232 327428 274238 327480
rect 267826 327292 267832 327344
rect 267884 327332 267890 327344
rect 268838 327332 268844 327344
rect 267884 327304 268844 327332
rect 267884 327292 267890 327304
rect 268838 327292 268844 327304
rect 268896 327292 268902 327344
rect 273438 327224 273444 327276
rect 273496 327264 273502 327276
rect 273898 327264 273904 327276
rect 273496 327236 273904 327264
rect 273496 327224 273502 327236
rect 273898 327224 273904 327236
rect 273956 327224 273962 327276
rect 336182 327196 336188 327208
rect 335832 327168 336188 327196
rect 335832 327140 335860 327168
rect 336182 327156 336188 327168
rect 336240 327156 336246 327208
rect 107470 327128 107476 327140
rect 107431 327100 107476 327128
rect 107470 327088 107476 327100
rect 107528 327088 107534 327140
rect 266814 327088 266820 327140
rect 266872 327128 266878 327140
rect 267458 327128 267464 327140
rect 266872 327100 267464 327128
rect 266872 327088 266878 327100
rect 267458 327088 267464 327100
rect 267516 327088 267522 327140
rect 272334 327088 272340 327140
rect 272392 327128 272398 327140
rect 272518 327128 272524 327140
rect 272392 327100 272524 327128
rect 272392 327088 272398 327100
rect 272518 327088 272524 327100
rect 272576 327088 272582 327140
rect 279510 327128 279516 327140
rect 279471 327100 279516 327128
rect 279510 327088 279516 327100
rect 279568 327088 279574 327140
rect 334526 327088 334532 327140
rect 334584 327128 334590 327140
rect 335170 327128 335176 327140
rect 334584 327100 335176 327128
rect 334584 327088 334590 327100
rect 335170 327088 335176 327100
rect 335228 327088 335234 327140
rect 335814 327088 335820 327140
rect 335872 327088 335878 327140
rect 257062 327060 257068 327072
rect 257023 327032 257068 327060
rect 257062 327020 257068 327032
rect 257120 327020 257126 327072
rect 295610 327060 295616 327072
rect 295571 327032 295616 327060
rect 295610 327020 295616 327032
rect 295668 327020 295674 327072
rect 341613 327063 341671 327069
rect 341613 327029 341625 327063
rect 341659 327060 341671 327063
rect 341702 327060 341708 327072
rect 341659 327032 341708 327060
rect 341659 327029 341671 327032
rect 341613 327023 341671 327029
rect 341702 327020 341708 327032
rect 341760 327020 341766 327072
rect 287422 326952 287428 327004
rect 287480 326992 287486 327004
rect 288066 326992 288072 327004
rect 287480 326964 288072 326992
rect 287480 326952 287486 326964
rect 288066 326952 288072 326964
rect 288124 326952 288130 327004
rect 270586 326680 270592 326732
rect 270644 326720 270650 326732
rect 271598 326720 271604 326732
rect 270644 326692 271604 326720
rect 270644 326680 270650 326692
rect 271598 326680 271604 326692
rect 271656 326680 271662 326732
rect 270770 326612 270776 326664
rect 270828 326652 270834 326664
rect 271414 326652 271420 326664
rect 270828 326624 271420 326652
rect 270828 326612 270834 326624
rect 271414 326612 271420 326624
rect 271472 326612 271478 326664
rect 297174 326544 297180 326596
rect 297232 326584 297238 326596
rect 297910 326584 297916 326596
rect 297232 326556 297916 326584
rect 297232 326544 297238 326556
rect 297910 326544 297916 326556
rect 297968 326544 297974 326596
rect 262398 326476 262404 326528
rect 262456 326516 262462 326528
rect 263318 326516 263324 326528
rect 262456 326488 263324 326516
rect 262456 326476 262462 326488
rect 263318 326476 263324 326488
rect 263376 326476 263382 326528
rect 282914 326476 282920 326528
rect 282972 326516 282978 326528
rect 284110 326516 284116 326528
rect 282972 326488 284116 326516
rect 282972 326476 282978 326488
rect 284110 326476 284116 326488
rect 284168 326476 284174 326528
rect 289906 326476 289912 326528
rect 289964 326516 289970 326528
rect 291102 326516 291108 326528
rect 289964 326488 291108 326516
rect 289964 326476 289970 326488
rect 291102 326476 291108 326488
rect 291160 326476 291166 326528
rect 291286 326476 291292 326528
rect 291344 326516 291350 326528
rect 292482 326516 292488 326528
rect 291344 326488 292488 326516
rect 291344 326476 291350 326488
rect 292482 326476 292488 326488
rect 292540 326476 292546 326528
rect 292758 326476 292764 326528
rect 292816 326516 292822 326528
rect 293770 326516 293776 326528
rect 292816 326488 293776 326516
rect 292816 326476 292822 326488
rect 293770 326476 293776 326488
rect 293828 326476 293834 326528
rect 297358 326476 297364 326528
rect 297416 326516 297422 326528
rect 298002 326516 298008 326528
rect 297416 326488 298008 326516
rect 297416 326476 297422 326488
rect 298002 326476 298008 326488
rect 298060 326476 298066 326528
rect 307846 326476 307852 326528
rect 307904 326516 307910 326528
rect 308950 326516 308956 326528
rect 307904 326488 308956 326516
rect 307904 326476 307910 326488
rect 308950 326476 308956 326488
rect 309008 326476 309014 326528
rect 311894 326476 311900 326528
rect 311952 326516 311958 326528
rect 313090 326516 313096 326528
rect 311952 326488 313096 326516
rect 311952 326476 311958 326488
rect 313090 326476 313096 326488
rect 313148 326476 313154 326528
rect 313274 326476 313280 326528
rect 313332 326516 313338 326528
rect 314562 326516 314568 326528
rect 313332 326488 314568 326516
rect 313332 326476 313338 326488
rect 314562 326476 314568 326488
rect 314620 326476 314626 326528
rect 315206 326476 315212 326528
rect 315264 326516 315270 326528
rect 315850 326516 315856 326528
rect 315264 326488 315856 326516
rect 315264 326476 315270 326488
rect 315850 326476 315856 326488
rect 315908 326476 315914 326528
rect 318794 326476 318800 326528
rect 318852 326516 318858 326528
rect 320082 326516 320088 326528
rect 318852 326488 320088 326516
rect 318852 326476 318858 326488
rect 320082 326476 320088 326488
rect 320140 326476 320146 326528
rect 259454 326408 259460 326460
rect 259512 326448 259518 326460
rect 260558 326448 260564 326460
rect 259512 326420 260564 326448
rect 259512 326408 259518 326420
rect 260558 326408 260564 326420
rect 260616 326408 260622 326460
rect 260834 326408 260840 326460
rect 260892 326448 260898 326460
rect 261846 326448 261852 326460
rect 260892 326420 261852 326448
rect 260892 326408 260898 326420
rect 261846 326408 261852 326420
rect 261904 326408 261910 326460
rect 262582 326408 262588 326460
rect 262640 326448 262646 326460
rect 263410 326448 263416 326460
rect 262640 326420 263416 326448
rect 262640 326408 262646 326420
rect 263410 326408 263416 326420
rect 263468 326408 263474 326460
rect 264974 326408 264980 326460
rect 265032 326448 265038 326460
rect 265894 326448 265900 326460
rect 265032 326420 265900 326448
rect 265032 326408 265038 326420
rect 265894 326408 265900 326420
rect 265952 326408 265958 326460
rect 266354 326408 266360 326460
rect 266412 326448 266418 326460
rect 267366 326448 267372 326460
rect 266412 326420 267372 326448
rect 266412 326408 266418 326420
rect 267366 326408 267372 326420
rect 267424 326408 267430 326460
rect 267734 326408 267740 326460
rect 267792 326448 267798 326460
rect 268930 326448 268936 326460
rect 267792 326420 268936 326448
rect 267792 326408 267798 326420
rect 268930 326408 268936 326420
rect 268988 326408 268994 326460
rect 269206 326408 269212 326460
rect 269264 326448 269270 326460
rect 270310 326448 270316 326460
rect 269264 326420 270316 326448
rect 269264 326408 269270 326420
rect 270310 326408 270316 326420
rect 270368 326408 270374 326460
rect 273438 326408 273444 326460
rect 273496 326448 273502 326460
rect 274266 326448 274272 326460
rect 273496 326420 274272 326448
rect 273496 326408 273502 326420
rect 274266 326408 274272 326420
rect 274324 326408 274330 326460
rect 275094 326408 275100 326460
rect 275152 326448 275158 326460
rect 275922 326448 275928 326460
rect 275152 326420 275928 326448
rect 275152 326408 275158 326420
rect 275922 326408 275928 326420
rect 275980 326408 275986 326460
rect 276290 326408 276296 326460
rect 276348 326448 276354 326460
rect 277026 326448 277032 326460
rect 276348 326420 277032 326448
rect 276348 326408 276354 326420
rect 277026 326408 277032 326420
rect 277084 326408 277090 326460
rect 277762 326408 277768 326460
rect 277820 326448 277826 326460
rect 278682 326448 278688 326460
rect 277820 326420 278688 326448
rect 277820 326408 277826 326420
rect 278682 326408 278688 326420
rect 278740 326408 278746 326460
rect 278774 326408 278780 326460
rect 278832 326448 278838 326460
rect 279878 326448 279884 326460
rect 278832 326420 279884 326448
rect 278832 326408 278838 326420
rect 279878 326408 279884 326420
rect 279936 326408 279942 326460
rect 280246 326408 280252 326460
rect 280304 326448 280310 326460
rect 281442 326448 281448 326460
rect 280304 326420 281448 326448
rect 280304 326408 280310 326420
rect 281442 326408 281448 326420
rect 281500 326408 281506 326460
rect 281626 326408 281632 326460
rect 281684 326448 281690 326460
rect 282546 326448 282552 326460
rect 281684 326420 282552 326448
rect 281684 326408 281690 326420
rect 282546 326408 282552 326420
rect 282604 326408 282610 326460
rect 283282 326408 283288 326460
rect 283340 326448 283346 326460
rect 284018 326448 284024 326460
rect 283340 326420 284024 326448
rect 283340 326408 283346 326420
rect 284018 326408 284024 326420
rect 284076 326408 284082 326460
rect 284386 326408 284392 326460
rect 284444 326448 284450 326460
rect 285582 326448 285588 326460
rect 284444 326420 285588 326448
rect 284444 326408 284450 326420
rect 285582 326408 285588 326420
rect 285640 326408 285646 326460
rect 285674 326408 285680 326460
rect 285732 326448 285738 326460
rect 286962 326448 286968 326460
rect 285732 326420 286968 326448
rect 285732 326408 285738 326420
rect 286962 326408 286968 326420
rect 287020 326408 287026 326460
rect 287698 326408 287704 326460
rect 287756 326448 287762 326460
rect 288342 326448 288348 326460
rect 287756 326420 288348 326448
rect 287756 326408 287762 326420
rect 288342 326408 288348 326420
rect 288400 326408 288406 326460
rect 288802 326408 288808 326460
rect 288860 326448 288866 326460
rect 289538 326448 289544 326460
rect 288860 326420 289544 326448
rect 288860 326408 288866 326420
rect 289538 326408 289544 326420
rect 289596 326408 289602 326460
rect 290090 326408 290096 326460
rect 290148 326448 290154 326460
rect 290918 326448 290924 326460
rect 290148 326420 290924 326448
rect 290148 326408 290154 326420
rect 290918 326408 290924 326420
rect 290976 326408 290982 326460
rect 291470 326408 291476 326460
rect 291528 326448 291534 326460
rect 292206 326448 292212 326460
rect 291528 326420 292212 326448
rect 291528 326408 291534 326420
rect 292206 326408 292212 326420
rect 292264 326408 292270 326460
rect 292942 326408 292948 326460
rect 293000 326448 293006 326460
rect 293586 326448 293592 326460
rect 293000 326420 293592 326448
rect 293000 326408 293006 326420
rect 293586 326408 293592 326420
rect 293644 326408 293650 326460
rect 294046 326408 294052 326460
rect 294104 326448 294110 326460
rect 295242 326448 295248 326460
rect 294104 326420 295248 326448
rect 294104 326408 294110 326420
rect 295242 326408 295248 326420
rect 295300 326408 295306 326460
rect 295886 326408 295892 326460
rect 295944 326448 295950 326460
rect 296530 326448 296536 326460
rect 295944 326420 296536 326448
rect 295944 326408 295950 326420
rect 296530 326408 296536 326420
rect 296588 326408 296594 326460
rect 298186 326408 298192 326460
rect 298244 326448 298250 326460
rect 299382 326448 299388 326460
rect 298244 326420 299388 326448
rect 298244 326408 298250 326420
rect 299382 326408 299388 326420
rect 299440 326408 299446 326460
rect 301222 326408 301228 326460
rect 301280 326448 301286 326460
rect 302142 326448 302148 326460
rect 301280 326420 302148 326448
rect 301280 326408 301286 326420
rect 302142 326408 302148 326420
rect 302200 326408 302206 326460
rect 302234 326408 302240 326460
rect 302292 326448 302298 326460
rect 303430 326448 303436 326460
rect 302292 326420 303436 326448
rect 302292 326408 302298 326420
rect 303430 326408 303436 326420
rect 303488 326408 303494 326460
rect 304074 326408 304080 326460
rect 304132 326448 304138 326460
rect 304810 326448 304816 326460
rect 304132 326420 304816 326448
rect 304132 326408 304138 326420
rect 304810 326408 304816 326420
rect 304868 326408 304874 326460
rect 305178 326408 305184 326460
rect 305236 326448 305242 326460
rect 306190 326448 306196 326460
rect 305236 326420 306196 326448
rect 305236 326408 305242 326420
rect 306190 326408 306196 326420
rect 306248 326408 306254 326460
rect 306466 326408 306472 326460
rect 306524 326448 306530 326460
rect 307662 326448 307668 326460
rect 306524 326420 307668 326448
rect 306524 326408 306530 326420
rect 307662 326408 307668 326420
rect 307720 326408 307726 326460
rect 308030 326408 308036 326460
rect 308088 326448 308094 326460
rect 308858 326448 308864 326460
rect 308088 326420 308864 326448
rect 308088 326408 308094 326420
rect 308858 326408 308864 326420
rect 308916 326408 308922 326460
rect 309134 326408 309140 326460
rect 309192 326448 309198 326460
rect 310238 326448 310244 326460
rect 309192 326420 310244 326448
rect 309192 326408 309198 326420
rect 310238 326408 310244 326420
rect 310296 326408 310302 326460
rect 311250 326408 311256 326460
rect 311308 326448 311314 326460
rect 311710 326448 311716 326460
rect 311308 326420 311716 326448
rect 311308 326408 311314 326420
rect 311710 326408 311716 326420
rect 311768 326408 311774 326460
rect 312078 326408 312084 326460
rect 312136 326448 312142 326460
rect 312814 326448 312820 326460
rect 312136 326420 312820 326448
rect 312136 326408 312142 326420
rect 312814 326408 312820 326420
rect 312872 326408 312878 326460
rect 313550 326408 313556 326460
rect 313608 326448 313614 326460
rect 314378 326448 314384 326460
rect 313608 326420 314384 326448
rect 313608 326408 313614 326420
rect 314378 326408 314384 326420
rect 314436 326408 314442 326460
rect 317966 326408 317972 326460
rect 318024 326448 318030 326460
rect 318426 326448 318432 326460
rect 318024 326420 318432 326448
rect 318024 326408 318030 326420
rect 318426 326408 318432 326420
rect 318484 326408 318490 326460
rect 319070 326408 319076 326460
rect 319128 326448 319134 326460
rect 319806 326448 319812 326460
rect 319128 326420 319812 326448
rect 319128 326408 319134 326420
rect 319806 326408 319812 326420
rect 319864 326408 319870 326460
rect 258718 326340 258724 326392
rect 258776 326380 258782 326392
rect 259270 326380 259276 326392
rect 258776 326352 259276 326380
rect 258776 326340 258782 326352
rect 259270 326340 259276 326352
rect 259328 326340 259334 326392
rect 259730 326340 259736 326392
rect 259788 326380 259794 326392
rect 260742 326380 260748 326392
rect 259788 326352 260748 326380
rect 259788 326340 259794 326352
rect 260742 326340 260748 326352
rect 260800 326340 260806 326392
rect 261202 326340 261208 326392
rect 261260 326380 261266 326392
rect 262030 326380 262036 326392
rect 261260 326352 262036 326380
rect 261260 326340 261266 326352
rect 262030 326340 262036 326352
rect 262088 326340 262094 326392
rect 262674 326340 262680 326392
rect 262732 326380 262738 326392
rect 263226 326380 263232 326392
rect 262732 326352 263232 326380
rect 262732 326340 262738 326352
rect 263226 326340 263232 326352
rect 263284 326340 263290 326392
rect 263594 326340 263600 326392
rect 263652 326380 263658 326392
rect 264790 326380 264796 326392
rect 263652 326352 264796 326380
rect 263652 326340 263658 326352
rect 264790 326340 264796 326352
rect 264848 326340 264854 326392
rect 265066 326340 265072 326392
rect 265124 326380 265130 326392
rect 265986 326380 265992 326392
rect 265124 326352 265992 326380
rect 265124 326340 265130 326352
rect 265986 326340 265992 326352
rect 266044 326340 266050 326392
rect 266630 326340 266636 326392
rect 266688 326380 266694 326392
rect 267550 326380 267556 326392
rect 266688 326352 267556 326380
rect 266688 326340 266694 326352
rect 267550 326340 267556 326352
rect 267608 326340 267614 326392
rect 268010 326340 268016 326392
rect 268068 326380 268074 326392
rect 268746 326380 268752 326392
rect 268068 326352 268752 326380
rect 268068 326340 268074 326352
rect 268746 326340 268752 326352
rect 268804 326340 268810 326392
rect 270678 326340 270684 326392
rect 270736 326380 270742 326392
rect 271782 326380 271788 326392
rect 270736 326352 271788 326380
rect 270736 326340 270742 326352
rect 271782 326340 271788 326352
rect 271840 326340 271846 326392
rect 271874 326340 271880 326392
rect 271932 326380 271938 326392
rect 272978 326380 272984 326392
rect 271932 326352 272984 326380
rect 271932 326340 271938 326352
rect 272978 326340 272984 326352
rect 273036 326340 273042 326392
rect 273714 326340 273720 326392
rect 273772 326380 273778 326392
rect 274358 326380 274364 326392
rect 273772 326352 274364 326380
rect 273772 326340 273778 326352
rect 274358 326340 274364 326352
rect 274416 326340 274422 326392
rect 274726 326340 274732 326392
rect 274784 326380 274790 326392
rect 275646 326380 275652 326392
rect 274784 326352 275652 326380
rect 274784 326340 274790 326352
rect 275646 326340 275652 326352
rect 275704 326340 275710 326392
rect 276658 326340 276664 326392
rect 276716 326380 276722 326392
rect 277210 326380 277216 326392
rect 276716 326352 277216 326380
rect 276716 326340 276722 326352
rect 277210 326340 277216 326352
rect 277268 326340 277274 326392
rect 277670 326340 277676 326392
rect 277728 326380 277734 326392
rect 278590 326380 278596 326392
rect 277728 326352 278596 326380
rect 277728 326340 277734 326352
rect 278590 326340 278596 326352
rect 278648 326340 278654 326392
rect 278866 326340 278872 326392
rect 278924 326380 278930 326392
rect 279786 326380 279792 326392
rect 278924 326352 279792 326380
rect 278924 326340 278930 326352
rect 279786 326340 279792 326352
rect 279844 326340 279850 326392
rect 280338 326340 280344 326392
rect 280396 326380 280402 326392
rect 281166 326380 281172 326392
rect 280396 326352 281172 326380
rect 280396 326340 280402 326352
rect 281166 326340 281172 326352
rect 281224 326340 281230 326392
rect 281718 326340 281724 326392
rect 281776 326380 281782 326392
rect 282454 326380 282460 326392
rect 281776 326352 282460 326380
rect 281776 326340 281782 326352
rect 282454 326340 282460 326352
rect 282512 326340 282518 326392
rect 283190 326340 283196 326392
rect 283248 326380 283254 326392
rect 283926 326380 283932 326392
rect 283248 326352 283932 326380
rect 283248 326340 283254 326352
rect 283926 326340 283932 326352
rect 283984 326340 283990 326392
rect 284294 326340 284300 326392
rect 284352 326380 284358 326392
rect 285490 326380 285496 326392
rect 284352 326352 285496 326380
rect 284352 326340 284358 326352
rect 285490 326340 285496 326352
rect 285548 326340 285554 326392
rect 285766 326340 285772 326392
rect 285824 326380 285830 326392
rect 286870 326380 286876 326392
rect 285824 326352 286876 326380
rect 285824 326340 285830 326352
rect 286870 326340 286876 326352
rect 286928 326340 286934 326392
rect 287606 326340 287612 326392
rect 287664 326380 287670 326392
rect 288158 326380 288164 326392
rect 287664 326352 288164 326380
rect 287664 326340 287670 326352
rect 288158 326340 288164 326352
rect 288216 326340 288222 326392
rect 288894 326340 288900 326392
rect 288952 326380 288958 326392
rect 289446 326380 289452 326392
rect 288952 326352 289452 326380
rect 288952 326340 288958 326352
rect 289446 326340 289452 326352
rect 289504 326340 289510 326392
rect 290182 326340 290188 326392
rect 290240 326380 290246 326392
rect 291010 326380 291016 326392
rect 290240 326352 291016 326380
rect 290240 326340 290246 326352
rect 291010 326340 291016 326352
rect 291068 326340 291074 326392
rect 291562 326340 291568 326392
rect 291620 326380 291626 326392
rect 292114 326380 292120 326392
rect 291620 326352 292120 326380
rect 291620 326340 291626 326352
rect 292114 326340 292120 326352
rect 292172 326340 292178 326392
rect 293034 326340 293040 326392
rect 293092 326380 293098 326392
rect 293494 326380 293500 326392
rect 293092 326352 293500 326380
rect 293092 326340 293098 326352
rect 293494 326340 293500 326352
rect 293552 326340 293558 326392
rect 294230 326340 294236 326392
rect 294288 326380 294294 326392
rect 295058 326380 295064 326392
rect 294288 326352 295064 326380
rect 294288 326340 294294 326352
rect 295058 326340 295064 326352
rect 295116 326340 295122 326392
rect 295334 326340 295340 326392
rect 295392 326380 295398 326392
rect 296622 326380 296628 326392
rect 295392 326352 296628 326380
rect 295392 326340 295398 326352
rect 296622 326340 296628 326352
rect 296680 326340 296686 326392
rect 296714 326340 296720 326392
rect 296772 326380 296778 326392
rect 297726 326380 297732 326392
rect 296772 326352 297732 326380
rect 296772 326340 296778 326352
rect 297726 326340 297732 326352
rect 297784 326340 297790 326392
rect 298370 326340 298376 326392
rect 298428 326380 298434 326392
rect 299290 326380 299296 326392
rect 298428 326352 299296 326380
rect 298428 326340 298434 326352
rect 299290 326340 299296 326352
rect 299348 326340 299354 326392
rect 302694 326340 302700 326392
rect 302752 326380 302758 326392
rect 303522 326380 303528 326392
rect 302752 326352 303528 326380
rect 302752 326340 302758 326352
rect 303522 326340 303528 326352
rect 303580 326340 303586 326392
rect 303798 326340 303804 326392
rect 303856 326380 303862 326392
rect 304626 326380 304632 326392
rect 303856 326352 304632 326380
rect 303856 326340 303862 326352
rect 304626 326340 304632 326352
rect 304684 326340 304690 326392
rect 305086 326340 305092 326392
rect 305144 326380 305150 326392
rect 306098 326380 306104 326392
rect 305144 326352 306104 326380
rect 305144 326340 305150 326352
rect 306098 326340 306104 326352
rect 306156 326340 306162 326392
rect 306558 326340 306564 326392
rect 306616 326380 306622 326392
rect 307478 326380 307484 326392
rect 306616 326352 307484 326380
rect 306616 326340 306622 326352
rect 307478 326340 307484 326352
rect 307536 326340 307542 326392
rect 308122 326340 308128 326392
rect 308180 326380 308186 326392
rect 308674 326380 308680 326392
rect 308180 326352 308680 326380
rect 308180 326340 308186 326352
rect 308674 326340 308680 326352
rect 308732 326340 308738 326392
rect 310606 326340 310612 326392
rect 310664 326380 310670 326392
rect 311802 326380 311808 326392
rect 310664 326352 311808 326380
rect 310664 326340 310670 326352
rect 311802 326340 311808 326352
rect 311860 326340 311866 326392
rect 312354 326340 312360 326392
rect 312412 326380 312418 326392
rect 312906 326380 312912 326392
rect 312412 326352 312912 326380
rect 312412 326340 312418 326352
rect 312906 326340 312912 326352
rect 312964 326340 312970 326392
rect 313642 326340 313648 326392
rect 313700 326380 313706 326392
rect 314286 326380 314292 326392
rect 313700 326352 314292 326380
rect 313700 326340 313706 326352
rect 314286 326340 314292 326352
rect 314344 326340 314350 326392
rect 314746 326340 314752 326392
rect 314804 326380 314810 326392
rect 315942 326380 315948 326392
rect 314804 326352 315948 326380
rect 314804 326340 314810 326352
rect 315942 326340 315948 326352
rect 316000 326340 316006 326392
rect 316218 326340 316224 326392
rect 316276 326380 316282 326392
rect 317230 326380 317236 326392
rect 316276 326352 317236 326380
rect 316276 326340 316282 326352
rect 317230 326340 317236 326352
rect 317288 326340 317294 326392
rect 318058 326340 318064 326392
rect 318116 326380 318122 326392
rect 318518 326380 318524 326392
rect 318116 326352 318524 326380
rect 318116 326340 318122 326352
rect 318518 326340 318524 326352
rect 318576 326340 318582 326392
rect 319162 326340 319168 326392
rect 319220 326380 319226 326392
rect 319714 326380 319720 326392
rect 319220 326352 319720 326380
rect 319220 326340 319226 326352
rect 319714 326340 319720 326352
rect 319772 326340 319778 326392
rect 320450 326340 320456 326392
rect 320508 326380 320514 326392
rect 321278 326380 321284 326392
rect 320508 326352 321284 326380
rect 320508 326340 320514 326352
rect 321278 326340 321284 326352
rect 321336 326340 321342 326392
rect 260926 326272 260932 326324
rect 260984 326312 260990 326324
rect 262122 326312 262128 326324
rect 260984 326284 262128 326312
rect 260984 326272 260990 326284
rect 262122 326272 262128 326284
rect 262180 326272 262186 326324
rect 262214 326272 262220 326324
rect 262272 326312 262278 326324
rect 263134 326312 263140 326324
rect 262272 326284 263140 326312
rect 262272 326272 262278 326284
rect 263134 326272 263140 326284
rect 263192 326272 263198 326324
rect 265158 326272 265164 326324
rect 265216 326312 265222 326324
rect 266170 326312 266176 326324
rect 265216 326284 266176 326312
rect 265216 326272 265222 326284
rect 266170 326272 266176 326284
rect 266228 326272 266234 326324
rect 266538 326272 266544 326324
rect 266596 326312 266602 326324
rect 267642 326312 267648 326324
rect 266596 326284 267648 326312
rect 266596 326272 266602 326284
rect 267642 326272 267648 326284
rect 267700 326272 267706 326324
rect 273254 326272 273260 326324
rect 273312 326312 273318 326324
rect 274542 326312 274548 326324
rect 273312 326284 274548 326312
rect 273312 326272 273318 326284
rect 274542 326272 274548 326284
rect 274600 326272 274606 326324
rect 276106 326272 276112 326324
rect 276164 326312 276170 326324
rect 276934 326312 276940 326324
rect 276164 326284 276940 326312
rect 276164 326272 276170 326284
rect 276934 326272 276940 326284
rect 276992 326272 276998 326324
rect 277394 326272 277400 326324
rect 277452 326312 277458 326324
rect 278314 326312 278320 326324
rect 277452 326284 278320 326312
rect 277452 326272 277458 326284
rect 278314 326272 278320 326284
rect 278372 326272 278378 326324
rect 279050 326272 279056 326324
rect 279108 326312 279114 326324
rect 280062 326312 280068 326324
rect 279108 326284 280068 326312
rect 279108 326272 279114 326284
rect 280062 326272 280068 326284
rect 280120 326272 280126 326324
rect 281534 326272 281540 326324
rect 281592 326312 281598 326324
rect 282730 326312 282736 326324
rect 281592 326284 282736 326312
rect 281592 326272 281598 326284
rect 282730 326272 282736 326284
rect 282788 326272 282794 326324
rect 283006 326272 283012 326324
rect 283064 326312 283070 326324
rect 284202 326312 284208 326324
rect 283064 326284 284208 326312
rect 283064 326272 283070 326284
rect 284202 326272 284208 326284
rect 284260 326272 284266 326324
rect 287330 326272 287336 326324
rect 287388 326312 287394 326324
rect 288250 326312 288256 326324
rect 287388 326284 288256 326312
rect 287388 326272 287394 326284
rect 288250 326272 288256 326284
rect 288308 326272 288314 326324
rect 288434 326272 288440 326324
rect 288492 326312 288498 326324
rect 289722 326312 289728 326324
rect 288492 326284 289728 326312
rect 288492 326272 288498 326284
rect 289722 326272 289728 326284
rect 289780 326272 289786 326324
rect 289814 326272 289820 326324
rect 289872 326312 289878 326324
rect 290826 326312 290832 326324
rect 289872 326284 290832 326312
rect 289872 326272 289878 326284
rect 290826 326272 290832 326284
rect 290884 326272 290890 326324
rect 291654 326272 291660 326324
rect 291712 326312 291718 326324
rect 292390 326312 292396 326324
rect 291712 326284 292396 326312
rect 291712 326272 291718 326284
rect 292390 326272 292396 326284
rect 292448 326272 292454 326324
rect 292850 326272 292856 326324
rect 292908 326312 292914 326324
rect 293678 326312 293684 326324
rect 292908 326284 293684 326312
rect 292908 326272 292914 326284
rect 293678 326272 293684 326284
rect 293736 326272 293742 326324
rect 303614 326272 303620 326324
rect 303672 326312 303678 326324
rect 304902 326312 304908 326324
rect 303672 326284 304908 326312
rect 303672 326272 303678 326284
rect 304902 326272 304908 326284
rect 304960 326272 304966 326324
rect 304994 326272 305000 326324
rect 305052 326312 305058 326324
rect 306282 326312 306288 326324
rect 305052 326284 306288 326312
rect 305052 326272 305058 326284
rect 306282 326272 306288 326284
rect 306340 326272 306346 326324
rect 307938 326272 307944 326324
rect 307996 326312 308002 326324
rect 308766 326312 308772 326324
rect 307996 326284 308772 326312
rect 307996 326272 308002 326284
rect 308766 326272 308772 326284
rect 308824 326272 308830 326324
rect 309226 326272 309232 326324
rect 309284 326312 309290 326324
rect 310422 326312 310428 326324
rect 309284 326284 310428 326312
rect 309284 326272 309290 326284
rect 310422 326272 310428 326284
rect 310480 326272 310486 326324
rect 312170 326272 312176 326324
rect 312228 326312 312234 326324
rect 312998 326312 313004 326324
rect 312228 326284 313004 326312
rect 312228 326272 312234 326284
rect 312998 326272 313004 326284
rect 313056 326272 313062 326324
rect 313366 326272 313372 326324
rect 313424 326312 313430 326324
rect 314470 326312 314476 326324
rect 313424 326284 314476 326312
rect 313424 326272 313430 326284
rect 314470 326272 314476 326284
rect 314528 326272 314534 326324
rect 317690 326272 317696 326324
rect 317748 326312 317754 326324
rect 318702 326312 318708 326324
rect 317748 326284 318708 326312
rect 317748 326272 317754 326284
rect 318702 326272 318708 326284
rect 318760 326272 318766 326324
rect 318978 326272 318984 326324
rect 319036 326312 319042 326324
rect 319990 326312 319996 326324
rect 319036 326284 319996 326312
rect 319036 326272 319042 326284
rect 319990 326272 319996 326284
rect 320048 326272 320054 326324
rect 256970 326204 256976 326256
rect 257028 326244 257034 326256
rect 257706 326244 257712 326256
rect 257028 326216 257712 326244
rect 257028 326204 257034 326216
rect 257706 326204 257712 326216
rect 257764 326204 257770 326256
rect 262490 326204 262496 326256
rect 262548 326244 262554 326256
rect 263502 326244 263508 326256
rect 262548 326216 263508 326244
rect 262548 326204 262554 326216
rect 263502 326204 263508 326216
rect 263560 326204 263566 326256
rect 292574 326204 292580 326256
rect 292632 326244 292638 326256
rect 293862 326244 293868 326256
rect 292632 326216 293868 326244
rect 292632 326204 292638 326216
rect 293862 326204 293868 326216
rect 293920 326204 293926 326256
rect 299658 326204 299664 326256
rect 299716 326244 299722 326256
rect 300486 326244 300492 326256
rect 299716 326216 300492 326244
rect 299716 326204 299722 326216
rect 300486 326204 300492 326216
rect 300544 326204 300550 326256
rect 300854 326204 300860 326256
rect 300912 326244 300918 326256
rect 301866 326244 301872 326256
rect 300912 326216 301872 326244
rect 300912 326204 300918 326216
rect 301866 326204 301872 326216
rect 301924 326204 301930 326256
rect 307754 326204 307760 326256
rect 307812 326244 307818 326256
rect 309042 326244 309048 326256
rect 307812 326216 309048 326244
rect 307812 326204 307818 326216
rect 309042 326204 309048 326216
rect 309100 326204 309106 326256
rect 310698 326204 310704 326256
rect 310756 326244 310762 326256
rect 311434 326244 311440 326256
rect 310756 326216 311440 326244
rect 310756 326204 310762 326216
rect 311434 326204 311440 326216
rect 311492 326204 311498 326256
rect 314838 326204 314844 326256
rect 314896 326244 314902 326256
rect 315574 326244 315580 326256
rect 314896 326216 315580 326244
rect 314896 326204 314902 326216
rect 315574 326204 315580 326216
rect 315632 326204 315638 326256
rect 256786 326136 256792 326188
rect 256844 326176 256850 326188
rect 257798 326176 257804 326188
rect 256844 326148 257804 326176
rect 256844 326136 256850 326148
rect 257798 326136 257804 326148
rect 257856 326136 257862 326188
rect 299474 326136 299480 326188
rect 299532 326176 299538 326188
rect 300394 326176 300400 326188
rect 299532 326148 300400 326176
rect 299532 326136 299538 326148
rect 300394 326136 300400 326148
rect 300452 326136 300458 326188
rect 299566 326068 299572 326120
rect 299624 326108 299630 326120
rect 300578 326108 300584 326120
rect 299624 326080 300584 326108
rect 299624 326068 299630 326080
rect 300578 326068 300584 326080
rect 300636 326068 300642 326120
rect 262769 325703 262827 325709
rect 262769 325669 262781 325703
rect 262815 325700 262827 325703
rect 262858 325700 262864 325712
rect 262815 325672 262864 325700
rect 262815 325669 262827 325672
rect 262769 325663 262827 325669
rect 262858 325660 262864 325672
rect 262916 325660 262922 325712
rect 318150 325660 318156 325712
rect 318208 325700 318214 325712
rect 318242 325700 318248 325712
rect 318208 325672 318248 325700
rect 318208 325660 318214 325672
rect 318242 325660 318248 325672
rect 318300 325660 318306 325712
rect 319438 325700 319444 325712
rect 319399 325672 319444 325700
rect 319438 325660 319444 325672
rect 319496 325660 319502 325712
rect 320266 325700 320272 325712
rect 320227 325672 320272 325700
rect 320266 325660 320272 325672
rect 320324 325660 320330 325712
rect 330754 325660 330760 325712
rect 330812 325700 330818 325712
rect 330938 325700 330944 325712
rect 330812 325672 330944 325700
rect 330812 325660 330818 325672
rect 330938 325660 330944 325672
rect 330996 325660 331002 325712
rect 335814 325632 335820 325644
rect 335775 325604 335820 325632
rect 335814 325592 335820 325604
rect 335872 325592 335878 325644
rect 296898 325524 296904 325576
rect 296956 325564 296962 325576
rect 297542 325564 297548 325576
rect 296956 325536 297548 325564
rect 296956 325524 296962 325536
rect 297542 325524 297548 325536
rect 297600 325524 297606 325576
rect 272242 324912 272248 324964
rect 272300 324952 272306 324964
rect 272794 324952 272800 324964
rect 272300 324924 272800 324952
rect 272300 324912 272306 324924
rect 272794 324912 272800 324924
rect 272852 324912 272858 324964
rect 268102 324708 268108 324760
rect 268160 324748 268166 324760
rect 268654 324748 268660 324760
rect 268160 324720 268660 324748
rect 268160 324708 268166 324720
rect 268654 324708 268660 324720
rect 268712 324708 268718 324760
rect 261110 324436 261116 324488
rect 261168 324476 261174 324488
rect 261570 324476 261576 324488
rect 261168 324448 261576 324476
rect 261168 324436 261174 324448
rect 261570 324436 261576 324448
rect 261628 324436 261634 324488
rect 2774 324164 2780 324216
rect 2832 324204 2838 324216
rect 4706 324204 4712 324216
rect 2832 324176 4712 324204
rect 2832 324164 2838 324176
rect 4706 324164 4712 324176
rect 4764 324164 4770 324216
rect 275002 323552 275008 323604
rect 275060 323592 275066 323604
rect 275554 323592 275560 323604
rect 275060 323564 275560 323592
rect 275060 323552 275066 323564
rect 275554 323552 275560 323564
rect 275612 323552 275618 323604
rect 298462 323552 298468 323604
rect 298520 323592 298526 323604
rect 299106 323592 299112 323604
rect 298520 323564 299112 323592
rect 298520 323552 298526 323564
rect 299106 323552 299112 323564
rect 299164 323552 299170 323604
rect 305454 323552 305460 323604
rect 305512 323592 305518 323604
rect 305914 323592 305920 323604
rect 305512 323564 305920 323592
rect 305512 323552 305518 323564
rect 305914 323552 305920 323564
rect 305972 323552 305978 323604
rect 309502 323552 309508 323604
rect 309560 323592 309566 323604
rect 310330 323592 310336 323604
rect 309560 323564 310336 323592
rect 309560 323552 309566 323564
rect 310330 323552 310336 323564
rect 310388 323552 310394 323604
rect 298094 323416 298100 323468
rect 298152 323456 298158 323468
rect 299014 323456 299020 323468
rect 298152 323428 299020 323456
rect 298152 323416 298158 323428
rect 299014 323416 299020 323428
rect 299072 323416 299078 323468
rect 262858 322192 262864 322244
rect 262916 322232 262922 322244
rect 263042 322232 263048 322244
rect 262916 322204 263048 322232
rect 262916 322192 262922 322204
rect 263042 322192 263048 322204
rect 263100 322192 263106 322244
rect 295613 322235 295671 322241
rect 295613 322201 295625 322235
rect 295659 322232 295671 322235
rect 296070 322232 296076 322244
rect 295659 322204 296076 322232
rect 295659 322201 295671 322204
rect 295613 322195 295671 322201
rect 296070 322192 296076 322204
rect 296128 322192 296134 322244
rect 244458 321580 244464 321632
rect 244516 321580 244522 321632
rect 244476 321496 244504 321580
rect 259730 321512 259736 321564
rect 259788 321552 259794 321564
rect 260374 321552 260380 321564
rect 259788 321524 260380 321552
rect 259788 321512 259794 321524
rect 260374 321512 260380 321524
rect 260432 321512 260438 321564
rect 309410 321512 309416 321564
rect 309468 321552 309474 321564
rect 310054 321552 310060 321564
rect 309468 321524 310060 321552
rect 309468 321512 309474 321524
rect 310054 321512 310060 321524
rect 310112 321512 310118 321564
rect 310882 321512 310888 321564
rect 310940 321552 310946 321564
rect 311342 321552 311348 321564
rect 310940 321524 311348 321552
rect 310940 321512 310946 321524
rect 311342 321512 311348 321524
rect 311400 321512 311406 321564
rect 244458 321444 244464 321496
rect 244516 321444 244522 321496
rect 266906 321444 266912 321496
rect 266964 321484 266970 321496
rect 267182 321484 267188 321496
rect 266964 321456 267188 321484
rect 266964 321444 266970 321456
rect 267182 321444 267188 321456
rect 267240 321444 267246 321496
rect 277578 321444 277584 321496
rect 277636 321484 277642 321496
rect 278222 321484 278228 321496
rect 277636 321456 278228 321484
rect 277636 321444 277642 321456
rect 278222 321444 278228 321456
rect 278280 321444 278286 321496
rect 302602 321444 302608 321496
rect 302660 321484 302666 321496
rect 303062 321484 303068 321496
rect 302660 321456 303068 321484
rect 302660 321444 302666 321456
rect 303062 321444 303068 321456
rect 303120 321444 303126 321496
rect 303890 321444 303896 321496
rect 303948 321484 303954 321496
rect 304442 321484 304448 321496
rect 303948 321456 304448 321484
rect 303948 321444 303954 321456
rect 304442 321444 304448 321456
rect 304500 321444 304506 321496
rect 100662 318832 100668 318844
rect 100623 318804 100668 318832
rect 100662 318792 100668 318804
rect 100720 318792 100726 318844
rect 231121 318835 231179 318841
rect 231121 318801 231133 318835
rect 231167 318832 231179 318835
rect 231210 318832 231216 318844
rect 231167 318804 231216 318832
rect 231167 318801 231179 318804
rect 231121 318795 231179 318801
rect 231210 318792 231216 318804
rect 231268 318792 231274 318844
rect 232314 318792 232320 318844
rect 232372 318832 232378 318844
rect 232406 318832 232412 318844
rect 232372 318804 232412 318832
rect 232372 318792 232378 318804
rect 232406 318792 232412 318804
rect 232464 318792 232470 318844
rect 232590 318792 232596 318844
rect 232648 318832 232654 318844
rect 232682 318832 232688 318844
rect 232648 318804 232688 318832
rect 232648 318792 232654 318804
rect 232682 318792 232688 318804
rect 232740 318792 232746 318844
rect 254673 318835 254731 318841
rect 254673 318801 254685 318835
rect 254719 318832 254731 318835
rect 254854 318832 254860 318844
rect 254719 318804 254860 318832
rect 254719 318801 254731 318804
rect 254673 318795 254731 318801
rect 254854 318792 254860 318804
rect 254912 318792 254918 318844
rect 265618 318792 265624 318844
rect 265676 318792 265682 318844
rect 272518 318792 272524 318844
rect 272576 318832 272582 318844
rect 272886 318832 272892 318844
rect 272576 318804 272892 318832
rect 272576 318792 272582 318804
rect 272886 318792 272892 318804
rect 272944 318792 272950 318844
rect 273806 318792 273812 318844
rect 273864 318832 273870 318844
rect 274082 318832 274088 318844
rect 273864 318804 274088 318832
rect 273864 318792 273870 318804
rect 274082 318792 274088 318804
rect 274140 318792 274146 318844
rect 280617 318835 280675 318841
rect 280617 318801 280629 318835
rect 280663 318832 280675 318835
rect 280982 318832 280988 318844
rect 280663 318804 280988 318832
rect 280663 318801 280675 318804
rect 280617 318795 280675 318801
rect 280982 318792 280988 318804
rect 281040 318792 281046 318844
rect 281905 318835 281963 318841
rect 281905 318801 281917 318835
rect 281951 318832 281963 318835
rect 282362 318832 282368 318844
rect 281951 318804 282368 318832
rect 281951 318801 281963 318804
rect 281905 318795 281963 318801
rect 282362 318792 282368 318804
rect 282420 318792 282426 318844
rect 344281 318835 344339 318841
rect 344281 318801 344293 318835
rect 344327 318832 344339 318835
rect 344370 318832 344376 318844
rect 344327 318804 344376 318832
rect 344327 318801 344339 318804
rect 344281 318795 344339 318801
rect 344370 318792 344376 318804
rect 344428 318792 344434 318844
rect 265636 318696 265664 318792
rect 315022 318724 315028 318776
rect 315080 318764 315086 318776
rect 315482 318764 315488 318776
rect 315080 318736 315488 318764
rect 315080 318724 315086 318736
rect 315482 318724 315488 318736
rect 315540 318724 315546 318776
rect 265802 318696 265808 318708
rect 265636 318668 265808 318696
rect 265802 318656 265808 318668
rect 265860 318656 265866 318708
rect 282638 318696 282644 318708
rect 282599 318668 282644 318696
rect 282638 318656 282644 318668
rect 282696 318656 282702 318708
rect 258718 317500 258724 317552
rect 258776 317540 258782 317552
rect 258902 317540 258908 317552
rect 258776 317512 258908 317540
rect 258776 317500 258782 317512
rect 258902 317500 258908 317512
rect 258960 317500 258966 317552
rect 257065 317475 257123 317481
rect 257065 317441 257077 317475
rect 257111 317472 257123 317475
rect 257154 317472 257160 317484
rect 257111 317444 257160 317472
rect 257111 317441 257123 317444
rect 257065 317435 257123 317441
rect 257154 317432 257160 317444
rect 257212 317432 257218 317484
rect 293310 317432 293316 317484
rect 293368 317472 293374 317484
rect 293402 317472 293408 317484
rect 293368 317444 293408 317472
rect 293368 317432 293374 317444
rect 293402 317432 293408 317444
rect 293460 317432 293466 317484
rect 293954 317432 293960 317484
rect 294012 317472 294018 317484
rect 294782 317472 294788 317484
rect 294012 317444 294788 317472
rect 294012 317432 294018 317444
rect 294782 317432 294788 317444
rect 294840 317432 294846 317484
rect 341610 317472 341616 317484
rect 341571 317444 341616 317472
rect 341610 317432 341616 317444
rect 341668 317432 341674 317484
rect 107470 317404 107476 317416
rect 107431 317376 107476 317404
rect 107470 317364 107476 317376
rect 107528 317364 107534 317416
rect 232314 317364 232320 317416
rect 232372 317404 232378 317416
rect 232406 317404 232412 317416
rect 232372 317376 232412 317404
rect 232372 317364 232378 317376
rect 232406 317364 232412 317376
rect 232464 317364 232470 317416
rect 244366 317404 244372 317416
rect 244327 317376 244372 317404
rect 244366 317364 244372 317376
rect 244424 317364 244430 317416
rect 260374 317404 260380 317416
rect 260335 317376 260380 317404
rect 260374 317364 260380 317376
rect 260432 317364 260438 317416
rect 261573 317407 261631 317413
rect 261573 317373 261585 317407
rect 261619 317404 261631 317407
rect 261662 317404 261668 317416
rect 261619 317376 261668 317404
rect 261619 317373 261631 317376
rect 261573 317367 261631 317373
rect 261662 317364 261668 317376
rect 261720 317364 261726 317416
rect 265802 317404 265808 317416
rect 265763 317376 265808 317404
rect 265802 317364 265808 317376
rect 265860 317364 265866 317416
rect 331766 317364 331772 317416
rect 331824 317404 331830 317416
rect 331858 317404 331864 317416
rect 331824 317376 331864 317404
rect 331824 317364 331830 317376
rect 331858 317364 331864 317376
rect 331916 317364 331922 317416
rect 333054 317364 333060 317416
rect 333112 317404 333118 317416
rect 333146 317404 333152 317416
rect 333112 317376 333152 317404
rect 333112 317364 333118 317376
rect 333146 317364 333152 317376
rect 333204 317364 333210 317416
rect 333238 317364 333244 317416
rect 333296 317404 333302 317416
rect 333330 317404 333336 317416
rect 333296 317376 333336 317404
rect 333296 317364 333302 317376
rect 333330 317364 333336 317376
rect 333388 317364 333394 317416
rect 339957 317407 340015 317413
rect 339957 317373 339969 317407
rect 340003 317404 340015 317407
rect 340138 317404 340144 317416
rect 340003 317376 340144 317404
rect 340003 317373 340015 317376
rect 339957 317367 340015 317373
rect 340138 317364 340144 317376
rect 340196 317364 340202 317416
rect 271966 316684 271972 316736
rect 272024 316724 272030 316736
rect 272702 316724 272708 316736
rect 272024 316696 272708 316724
rect 272024 316684 272030 316696
rect 272702 316684 272708 316696
rect 272760 316684 272766 316736
rect 284570 316548 284576 316600
rect 284628 316548 284634 316600
rect 316126 316548 316132 316600
rect 316184 316588 316190 316600
rect 316862 316588 316868 316600
rect 316184 316560 316868 316588
rect 316184 316548 316190 316560
rect 316862 316548 316868 316560
rect 316920 316548 316926 316600
rect 284588 316520 284616 316548
rect 285030 316520 285036 316532
rect 284588 316492 285036 316520
rect 285030 316480 285036 316492
rect 285088 316480 285094 316532
rect 319438 316072 319444 316124
rect 319496 316112 319502 316124
rect 319622 316112 319628 316124
rect 319496 316084 319628 316112
rect 319496 316072 319502 316084
rect 319622 316072 319628 316084
rect 319680 316072 319686 316124
rect 301038 316004 301044 316056
rect 301096 316044 301102 316056
rect 301774 316044 301780 316056
rect 301096 316016 301780 316044
rect 301096 316004 301102 316016
rect 301774 316004 301780 316016
rect 301832 316004 301838 316056
rect 330570 316004 330576 316056
rect 330628 316044 330634 316056
rect 330754 316044 330760 316056
rect 330628 316016 330760 316044
rect 330628 316004 330634 316016
rect 330754 316004 330760 316016
rect 330812 316004 330818 316056
rect 335817 316047 335875 316053
rect 335817 316013 335829 316047
rect 335863 316044 335875 316047
rect 335998 316044 336004 316056
rect 335863 316016 336004 316044
rect 335863 316013 335875 316016
rect 335817 316007 335875 316013
rect 335998 316004 336004 316016
rect 336056 316004 336062 316056
rect 258813 315979 258871 315985
rect 258813 315945 258825 315979
rect 258859 315976 258871 315979
rect 258902 315976 258908 315988
rect 258859 315948 258908 315976
rect 258859 315945 258871 315948
rect 258813 315939 258871 315945
rect 258902 315936 258908 315948
rect 258960 315936 258966 315988
rect 319438 315976 319444 315988
rect 319399 315948 319444 315976
rect 319438 315936 319444 315948
rect 319496 315936 319502 315988
rect 320266 315976 320272 315988
rect 320227 315948 320272 315976
rect 320266 315936 320272 315948
rect 320324 315936 320330 315988
rect 317874 315188 317880 315240
rect 317932 315228 317938 315240
rect 318242 315228 318248 315240
rect 317932 315200 318248 315228
rect 317932 315188 317938 315200
rect 318242 315188 318248 315200
rect 318300 315188 318306 315240
rect 285858 313896 285864 313948
rect 285916 313936 285922 313948
rect 286502 313936 286508 313948
rect 285916 313908 286508 313936
rect 285916 313896 285922 313908
rect 286502 313896 286508 313908
rect 286560 313896 286566 313948
rect 263778 313488 263784 313540
rect 263836 313528 263842 313540
rect 264514 313528 264520 313540
rect 263836 313500 264520 313528
rect 263836 313488 263842 313500
rect 264514 313488 264520 313500
rect 264572 313488 264578 313540
rect 322290 312672 322296 312724
rect 322348 312712 322354 312724
rect 322566 312712 322572 312724
rect 322348 312684 322572 312712
rect 322348 312672 322354 312684
rect 322566 312672 322572 312684
rect 322624 312672 322630 312724
rect 231210 311924 231216 311976
rect 231268 311924 231274 311976
rect 289262 311964 289268 311976
rect 289188 311936 289268 311964
rect 231228 311772 231256 311924
rect 289188 311840 289216 311936
rect 289262 311924 289268 311936
rect 289320 311924 289326 311976
rect 344186 311856 344192 311908
rect 344244 311896 344250 311908
rect 344370 311896 344376 311908
rect 344244 311868 344376 311896
rect 344244 311856 344250 311868
rect 344370 311856 344376 311868
rect 344428 311856 344434 311908
rect 289170 311788 289176 311840
rect 289228 311788 289234 311840
rect 231210 311720 231216 311772
rect 231268 311720 231274 311772
rect 244366 311488 244372 311500
rect 244327 311460 244372 311488
rect 244366 311448 244372 311460
rect 244424 311448 244430 311500
rect 322290 311108 322296 311160
rect 322348 311148 322354 311160
rect 322566 311148 322572 311160
rect 322348 311120 322572 311148
rect 322348 311108 322354 311120
rect 322566 311108 322572 311120
rect 322624 311108 322630 311160
rect 310054 309884 310060 309936
rect 310112 309884 310118 309936
rect 311342 309884 311348 309936
rect 311400 309884 311406 309936
rect 310072 309800 310100 309884
rect 311360 309800 311388 309884
rect 310054 309748 310060 309800
rect 310112 309748 310118 309800
rect 311342 309748 311348 309800
rect 311400 309748 311406 309800
rect 280890 309136 280896 309188
rect 280948 309176 280954 309188
rect 280982 309176 280988 309188
rect 280948 309148 280988 309176
rect 280948 309136 280954 309148
rect 280982 309136 280988 309148
rect 281040 309136 281046 309188
rect 282638 309176 282644 309188
rect 282599 309148 282644 309176
rect 282638 309136 282644 309148
rect 282696 309136 282702 309188
rect 293310 309136 293316 309188
rect 293368 309176 293374 309188
rect 293405 309179 293463 309185
rect 293405 309176 293417 309179
rect 293368 309148 293417 309176
rect 293368 309136 293374 309148
rect 293405 309145 293417 309148
rect 293451 309145 293463 309179
rect 293405 309139 293463 309145
rect 100662 309108 100668 309120
rect 100623 309080 100668 309108
rect 100662 309068 100668 309080
rect 100720 309068 100726 309120
rect 238018 309108 238024 309120
rect 237979 309080 238024 309108
rect 238018 309068 238024 309080
rect 238076 309068 238082 309120
rect 246390 309068 246396 309120
rect 246448 309068 246454 309120
rect 253106 309068 253112 309120
rect 253164 309108 253170 309120
rect 253198 309108 253204 309120
rect 253164 309080 253204 309108
rect 253164 309068 253170 309080
rect 253198 309068 253204 309080
rect 253256 309068 253262 309120
rect 254670 309068 254676 309120
rect 254728 309108 254734 309120
rect 254854 309108 254860 309120
rect 254728 309080 254860 309108
rect 254728 309068 254734 309080
rect 254854 309068 254860 309080
rect 254912 309068 254918 309120
rect 257062 309068 257068 309120
rect 257120 309108 257126 309120
rect 257154 309108 257160 309120
rect 257120 309080 257160 309108
rect 257120 309068 257126 309080
rect 257154 309068 257160 309080
rect 257212 309068 257218 309120
rect 326246 309068 326252 309120
rect 326304 309108 326310 309120
rect 326338 309108 326344 309120
rect 326304 309080 326344 309108
rect 326304 309068 326310 309080
rect 326338 309068 326344 309080
rect 326396 309068 326402 309120
rect 246408 309040 246436 309068
rect 246482 309040 246488 309052
rect 246408 309012 246488 309040
rect 246482 309000 246488 309012
rect 246540 309000 246546 309052
rect 265802 307884 265808 307896
rect 265763 307856 265808 307884
rect 265802 307844 265808 307856
rect 265860 307844 265866 307896
rect 107470 307816 107476 307828
rect 107431 307788 107476 307816
rect 107470 307776 107476 307788
rect 107528 307776 107534 307828
rect 260374 307816 260380 307828
rect 260335 307788 260380 307816
rect 260374 307776 260380 307788
rect 260432 307776 260438 307828
rect 329006 307776 329012 307828
rect 329064 307816 329070 307828
rect 329098 307816 329104 307828
rect 329064 307788 329104 307816
rect 329064 307776 329070 307788
rect 329098 307776 329104 307788
rect 329156 307776 329162 307828
rect 339954 307816 339960 307828
rect 339915 307788 339960 307816
rect 339954 307776 339960 307788
rect 340012 307776 340018 307828
rect 264514 307748 264520 307760
rect 264475 307720 264520 307748
rect 264514 307708 264520 307720
rect 264572 307708 264578 307760
rect 265802 307748 265808 307760
rect 265763 307720 265808 307748
rect 265802 307708 265808 307720
rect 265860 307708 265866 307760
rect 316862 307748 316868 307760
rect 316823 307720 316868 307748
rect 316862 307708 316868 307720
rect 316920 307708 316926 307760
rect 318058 307028 318064 307080
rect 318116 307068 318122 307080
rect 318334 307068 318340 307080
rect 318116 307040 318340 307068
rect 318116 307028 318122 307040
rect 318334 307028 318340 307040
rect 318392 307028 318398 307080
rect 293402 306388 293408 306400
rect 293363 306360 293408 306388
rect 293402 306348 293408 306360
rect 293460 306348 293466 306400
rect 319441 306391 319499 306397
rect 319441 306357 319453 306391
rect 319487 306388 319499 306391
rect 319622 306388 319628 306400
rect 319487 306360 319628 306388
rect 319487 306357 319499 306360
rect 319441 306351 319499 306357
rect 319622 306348 319628 306360
rect 319680 306348 319686 306400
rect 320269 306391 320327 306397
rect 320269 306357 320281 306391
rect 320315 306388 320327 306391
rect 321094 306388 321100 306400
rect 320315 306360 321100 306388
rect 320315 306357 320327 306360
rect 320269 306351 320327 306357
rect 321094 306348 321100 306360
rect 321152 306348 321158 306400
rect 335814 306348 335820 306400
rect 335872 306388 335878 306400
rect 335998 306388 336004 306400
rect 335872 306360 336004 306388
rect 335872 306348 335878 306360
rect 335998 306348 336004 306360
rect 336056 306348 336062 306400
rect 267182 304308 267188 304360
rect 267240 304308 267246 304360
rect 268654 304308 268660 304360
rect 268712 304308 268718 304360
rect 267200 304224 267228 304308
rect 268672 304224 268700 304308
rect 267182 304172 267188 304224
rect 267240 304172 267246 304224
rect 268654 304172 268660 304224
rect 268712 304172 268718 304224
rect 257062 302920 257068 302932
rect 257023 302892 257068 302920
rect 257062 302880 257068 302892
rect 257120 302880 257126 302932
rect 341610 302200 341616 302252
rect 341668 302200 341674 302252
rect 341628 302104 341656 302200
rect 341702 302104 341708 302116
rect 341628 302076 341708 302104
rect 341702 302064 341708 302076
rect 341760 302064 341766 302116
rect 100662 299520 100668 299532
rect 100623 299492 100668 299520
rect 100662 299480 100668 299492
rect 100720 299480 100726 299532
rect 238018 299520 238024 299532
rect 237979 299492 238024 299520
rect 238018 299480 238024 299492
rect 238076 299480 238082 299532
rect 244918 299480 244924 299532
rect 244976 299520 244982 299532
rect 245010 299520 245016 299532
rect 244976 299492 245016 299520
rect 244976 299480 244982 299492
rect 245010 299480 245016 299492
rect 245068 299480 245074 299532
rect 254670 299480 254676 299532
rect 254728 299480 254734 299532
rect 261570 299520 261576 299532
rect 261531 299492 261576 299520
rect 261570 299480 261576 299492
rect 261628 299480 261634 299532
rect 322198 299480 322204 299532
rect 322256 299520 322262 299532
rect 322290 299520 322296 299532
rect 322256 299492 322296 299520
rect 322256 299480 322262 299492
rect 322290 299480 322296 299492
rect 322348 299480 322354 299532
rect 231210 299452 231216 299464
rect 231171 299424 231216 299452
rect 231210 299412 231216 299424
rect 231268 299412 231274 299464
rect 231946 299412 231952 299464
rect 232004 299452 232010 299464
rect 232038 299452 232044 299464
rect 232004 299424 232044 299452
rect 232004 299412 232010 299424
rect 232038 299412 232044 299424
rect 232096 299412 232102 299464
rect 232314 299412 232320 299464
rect 232372 299452 232378 299464
rect 232406 299452 232412 299464
rect 232372 299424 232412 299452
rect 232372 299412 232378 299424
rect 232406 299412 232412 299424
rect 232464 299412 232470 299464
rect 240686 299452 240692 299464
rect 240647 299424 240692 299452
rect 240686 299412 240692 299424
rect 240744 299412 240750 299464
rect 246390 299412 246396 299464
rect 246448 299452 246454 299464
rect 246482 299452 246488 299464
rect 246448 299424 246488 299452
rect 246448 299412 246454 299424
rect 246482 299412 246488 299424
rect 246540 299412 246546 299464
rect 254688 299384 254716 299480
rect 260282 299452 260288 299464
rect 260243 299424 260288 299452
rect 260282 299412 260288 299424
rect 260340 299412 260346 299464
rect 331766 299412 331772 299464
rect 331824 299452 331830 299464
rect 331858 299452 331864 299464
rect 331824 299424 331864 299452
rect 331824 299412 331830 299424
rect 331858 299412 331864 299424
rect 331916 299412 331922 299464
rect 333238 299412 333244 299464
rect 333296 299452 333302 299464
rect 333330 299452 333336 299464
rect 333296 299424 333336 299452
rect 333296 299412 333302 299424
rect 333330 299412 333336 299424
rect 333388 299412 333394 299464
rect 334526 299412 334532 299464
rect 334584 299452 334590 299464
rect 334618 299452 334624 299464
rect 334584 299424 334624 299452
rect 334584 299412 334590 299424
rect 334618 299412 334624 299424
rect 334676 299412 334682 299464
rect 339954 299412 339960 299464
rect 340012 299452 340018 299464
rect 340138 299452 340144 299464
rect 340012 299424 340144 299452
rect 340012 299412 340018 299424
rect 340138 299412 340144 299424
rect 340196 299412 340202 299464
rect 341702 299412 341708 299464
rect 341760 299412 341766 299464
rect 345382 299412 345388 299464
rect 345440 299412 345446 299464
rect 254854 299384 254860 299396
rect 254688 299356 254860 299384
rect 254854 299344 254860 299356
rect 254912 299344 254918 299396
rect 341720 299328 341748 299412
rect 345400 299328 345428 299412
rect 341702 299276 341708 299328
rect 341760 299276 341766 299328
rect 345382 299276 345388 299328
rect 345440 299276 345446 299328
rect 258810 298120 258816 298172
rect 258868 298160 258874 298172
rect 258868 298132 258913 298160
rect 258868 298120 258874 298132
rect 264514 298120 264520 298172
rect 264572 298160 264578 298172
rect 264572 298132 264617 298160
rect 264572 298120 264578 298132
rect 265802 298120 265808 298172
rect 265860 298160 265866 298172
rect 265860 298132 265905 298160
rect 265860 298120 265866 298132
rect 293310 298120 293316 298172
rect 293368 298160 293374 298172
rect 293402 298160 293408 298172
rect 293368 298132 293408 298160
rect 293368 298120 293374 298132
rect 293402 298120 293408 298132
rect 293460 298120 293466 298172
rect 316865 298163 316923 298169
rect 316865 298129 316877 298163
rect 316911 298160 316923 298163
rect 316954 298160 316960 298172
rect 316911 298132 316960 298160
rect 316911 298129 316923 298132
rect 316865 298123 316923 298129
rect 316954 298120 316960 298132
rect 317012 298120 317018 298172
rect 107470 298092 107476 298104
rect 107431 298064 107476 298092
rect 107470 298052 107476 298064
rect 107528 298052 107534 298104
rect 231946 298052 231952 298104
rect 232004 298092 232010 298104
rect 232038 298092 232044 298104
rect 232004 298064 232044 298092
rect 232004 298052 232010 298064
rect 232038 298052 232044 298064
rect 232096 298052 232102 298104
rect 232406 298092 232412 298104
rect 232367 298064 232412 298092
rect 232406 298052 232412 298064
rect 232464 298052 232470 298104
rect 245010 298092 245016 298104
rect 244971 298064 245016 298092
rect 245010 298052 245016 298064
rect 245068 298052 245074 298104
rect 319622 298092 319628 298104
rect 319583 298064 319628 298092
rect 319622 298052 319628 298064
rect 319680 298052 319686 298104
rect 321094 298092 321100 298104
rect 321055 298064 321100 298092
rect 321094 298052 321100 298064
rect 321152 298052 321158 298104
rect 333238 298052 333244 298104
rect 333296 298092 333302 298104
rect 333330 298092 333336 298104
rect 333296 298064 333336 298092
rect 333296 298052 333302 298064
rect 333330 298052 333336 298064
rect 333388 298052 333394 298104
rect 339954 298092 339960 298104
rect 339915 298064 339960 298092
rect 339954 298052 339960 298064
rect 340012 298052 340018 298104
rect 335906 296692 335912 296744
rect 335964 296732 335970 296744
rect 335998 296732 336004 296744
rect 335964 296704 336004 296732
rect 335964 296692 335970 296704
rect 335998 296692 336004 296704
rect 336056 296692 336062 296744
rect 257065 294491 257123 294497
rect 257065 294457 257077 294491
rect 257111 294488 257123 294491
rect 257154 294488 257160 294500
rect 257111 294460 257160 294488
rect 257111 294457 257123 294460
rect 257065 294451 257123 294457
rect 257154 294448 257160 294460
rect 257212 294448 257218 294500
rect 232682 292612 232688 292664
rect 232740 292612 232746 292664
rect 232700 292528 232728 292612
rect 232682 292476 232688 292528
rect 232740 292476 232746 292528
rect 333146 290000 333152 290012
rect 333107 289972 333152 290000
rect 333146 289960 333152 289972
rect 333204 289960 333210 290012
rect 231210 289864 231216 289876
rect 231171 289836 231216 289864
rect 231210 289824 231216 289836
rect 231268 289824 231274 289876
rect 240686 289864 240692 289876
rect 240647 289836 240692 289864
rect 240686 289824 240692 289836
rect 240744 289824 240750 289876
rect 244366 289824 244372 289876
rect 244424 289864 244430 289876
rect 244458 289864 244464 289876
rect 244424 289836 244464 289864
rect 244424 289824 244430 289836
rect 244458 289824 244464 289836
rect 244516 289824 244522 289876
rect 253014 289824 253020 289876
rect 253072 289864 253078 289876
rect 253198 289864 253204 289876
rect 253072 289836 253204 289864
rect 253072 289824 253078 289836
rect 253198 289824 253204 289836
rect 253256 289824 253262 289876
rect 260285 289867 260343 289873
rect 260285 289833 260297 289867
rect 260331 289864 260343 289867
rect 260374 289864 260380 289876
rect 260331 289836 260380 289864
rect 260331 289833 260343 289836
rect 260285 289827 260343 289833
rect 260374 289824 260380 289836
rect 260432 289824 260438 289876
rect 322198 289824 322204 289876
rect 322256 289824 322262 289876
rect 331858 289864 331864 289876
rect 331784 289836 331864 289864
rect 100662 289796 100668 289808
rect 100623 289768 100668 289796
rect 100662 289756 100668 289768
rect 100720 289756 100726 289808
rect 238018 289796 238024 289808
rect 237979 289768 238024 289796
rect 238018 289756 238024 289768
rect 238076 289756 238082 289808
rect 261478 289756 261484 289808
rect 261536 289796 261542 289808
rect 261570 289796 261576 289808
rect 261536 289768 261576 289796
rect 261536 289756 261542 289768
rect 261570 289756 261576 289768
rect 261628 289756 261634 289808
rect 322216 289740 322244 289824
rect 331784 289808 331812 289836
rect 331858 289824 331864 289836
rect 331916 289824 331922 289876
rect 334618 289864 334624 289876
rect 334544 289836 334624 289864
rect 334544 289808 334572 289836
rect 334618 289824 334624 289836
rect 334676 289824 334682 289876
rect 331766 289756 331772 289808
rect 331824 289756 331830 289808
rect 334526 289756 334532 289808
rect 334584 289756 334590 289808
rect 322198 289688 322204 289740
rect 322256 289688 322262 289740
rect 321094 288504 321100 288516
rect 321055 288476 321100 288504
rect 321094 288464 321100 288476
rect 321152 288464 321158 288516
rect 329006 288464 329012 288516
rect 329064 288504 329070 288516
rect 329190 288504 329196 288516
rect 329064 288476 329196 288504
rect 329064 288464 329070 288476
rect 329190 288464 329196 288476
rect 329248 288464 329254 288516
rect 330570 288504 330576 288516
rect 330496 288476 330576 288504
rect 330496 288448 330524 288476
rect 330570 288464 330576 288476
rect 330628 288464 330634 288516
rect 335814 288464 335820 288516
rect 335872 288504 335878 288516
rect 335998 288504 336004 288516
rect 335872 288476 336004 288504
rect 335872 288464 335878 288476
rect 335998 288464 336004 288476
rect 336056 288464 336062 288516
rect 107470 288436 107476 288448
rect 107431 288408 107476 288436
rect 107470 288396 107476 288408
rect 107528 288396 107534 288448
rect 232406 288436 232412 288448
rect 232367 288408 232412 288436
rect 232406 288396 232412 288408
rect 232464 288396 232470 288448
rect 254854 288396 254860 288448
rect 254912 288436 254918 288448
rect 254946 288436 254952 288448
rect 254912 288408 254952 288436
rect 254912 288396 254918 288408
rect 254946 288396 254952 288408
rect 255004 288396 255010 288448
rect 293218 288396 293224 288448
rect 293276 288436 293282 288448
rect 293310 288436 293316 288448
rect 293276 288408 293316 288436
rect 293276 288396 293282 288408
rect 293310 288396 293316 288408
rect 293368 288396 293374 288448
rect 330478 288396 330484 288448
rect 330536 288396 330542 288448
rect 333146 288436 333152 288448
rect 333107 288408 333152 288436
rect 333146 288396 333152 288408
rect 333204 288396 333210 288448
rect 246390 288368 246396 288380
rect 246351 288340 246396 288368
rect 246390 288328 246396 288340
rect 246448 288328 246454 288380
rect 265802 288368 265808 288380
rect 265763 288340 265808 288368
rect 265802 288328 265808 288340
rect 265860 288328 265866 288380
rect 319622 287076 319628 287088
rect 319583 287048 319628 287076
rect 319622 287036 319628 287048
rect 319680 287036 319686 287088
rect 326246 287036 326252 287088
rect 326304 287076 326310 287088
rect 326430 287076 326436 287088
rect 326304 287048 326436 287076
rect 326304 287036 326310 287048
rect 326430 287036 326436 287048
rect 326488 287036 326494 287088
rect 258721 287011 258779 287017
rect 258721 286977 258733 287011
rect 258767 287008 258779 287011
rect 258902 287008 258908 287020
rect 258767 286980 258908 287008
rect 258767 286977 258779 286980
rect 258721 286971 258779 286977
rect 258902 286968 258908 286980
rect 258960 286968 258966 287020
rect 339957 282863 340015 282869
rect 339957 282829 339969 282863
rect 340003 282860 340015 282863
rect 340046 282860 340052 282872
rect 340003 282832 340052 282860
rect 340003 282829 340015 282832
rect 339957 282823 340015 282829
rect 340046 282820 340052 282832
rect 340104 282820 340110 282872
rect 100662 280208 100668 280220
rect 100623 280180 100668 280208
rect 100662 280168 100668 280180
rect 100720 280168 100726 280220
rect 238018 280208 238024 280220
rect 237979 280180 238024 280208
rect 238018 280168 238024 280180
rect 238076 280168 238082 280220
rect 254762 280168 254768 280220
rect 254820 280208 254826 280220
rect 254854 280208 254860 280220
rect 254820 280180 254860 280208
rect 254820 280168 254826 280180
rect 254854 280168 254860 280180
rect 254912 280168 254918 280220
rect 2774 280100 2780 280152
rect 2832 280140 2838 280152
rect 5442 280140 5448 280152
rect 2832 280112 5448 280140
rect 2832 280100 2838 280112
rect 5442 280100 5448 280112
rect 5500 280100 5506 280152
rect 231210 280140 231216 280152
rect 231171 280112 231216 280140
rect 231210 280100 231216 280112
rect 231268 280100 231274 280152
rect 232038 280100 232044 280152
rect 232096 280140 232102 280152
rect 232130 280140 232136 280152
rect 232096 280112 232136 280140
rect 232096 280100 232102 280112
rect 232130 280100 232136 280112
rect 232188 280100 232194 280152
rect 240686 280140 240692 280152
rect 240647 280112 240692 280140
rect 240686 280100 240692 280112
rect 240744 280100 240750 280152
rect 246022 280140 246028 280152
rect 245983 280112 246028 280140
rect 246022 280100 246028 280112
rect 246080 280100 246086 280152
rect 257154 280140 257160 280152
rect 257115 280112 257160 280140
rect 257154 280100 257160 280112
rect 257212 280100 257218 280152
rect 330478 280100 330484 280152
rect 330536 280140 330542 280152
rect 330570 280140 330576 280152
rect 330536 280112 330576 280140
rect 330536 280100 330542 280112
rect 330570 280100 330576 280112
rect 330628 280100 330634 280152
rect 331766 280100 331772 280152
rect 331824 280140 331830 280152
rect 331858 280140 331864 280152
rect 331824 280112 331864 280140
rect 331824 280100 331830 280112
rect 331858 280100 331864 280112
rect 331916 280100 331922 280152
rect 333238 280100 333244 280152
rect 333296 280140 333302 280152
rect 333330 280140 333336 280152
rect 333296 280112 333336 280140
rect 333296 280100 333302 280112
rect 333330 280100 333336 280112
rect 333388 280100 333394 280152
rect 334526 280100 334532 280152
rect 334584 280140 334590 280152
rect 334618 280140 334624 280152
rect 334584 280112 334624 280140
rect 334584 280100 334590 280112
rect 334618 280100 334624 280112
rect 334676 280100 334682 280152
rect 340046 280100 340052 280152
rect 340104 280140 340110 280152
rect 340138 280140 340144 280152
rect 340104 280112 340144 280140
rect 340104 280100 340110 280112
rect 340138 280100 340144 280112
rect 340196 280100 340202 280152
rect 265802 278848 265808 278860
rect 265763 278820 265808 278848
rect 265802 278808 265808 278820
rect 265860 278808 265866 278860
rect 244458 278740 244464 278792
rect 244516 278780 244522 278792
rect 244642 278780 244648 278792
rect 244516 278752 244648 278780
rect 244516 278740 244522 278752
rect 244642 278740 244648 278752
rect 244700 278740 244706 278792
rect 244918 278740 244924 278792
rect 244976 278780 244982 278792
rect 245013 278783 245071 278789
rect 245013 278780 245025 278783
rect 244976 278752 245025 278780
rect 244976 278740 244982 278752
rect 245013 278749 245025 278752
rect 245059 278749 245071 278783
rect 245013 278743 245071 278749
rect 246393 278783 246451 278789
rect 246393 278749 246405 278783
rect 246439 278780 246451 278783
rect 246482 278780 246488 278792
rect 246439 278752 246488 278780
rect 246439 278749 246451 278752
rect 246393 278743 246451 278749
rect 246482 278740 246488 278752
rect 246540 278740 246546 278792
rect 257154 278780 257160 278792
rect 257115 278752 257160 278780
rect 257154 278740 257160 278752
rect 257212 278740 257218 278792
rect 293126 278740 293132 278792
rect 293184 278780 293190 278792
rect 293310 278780 293316 278792
rect 293184 278752 293316 278780
rect 293184 278740 293190 278752
rect 293310 278740 293316 278752
rect 293368 278740 293374 278792
rect 329006 278740 329012 278792
rect 329064 278780 329070 278792
rect 329190 278780 329196 278792
rect 329064 278752 329196 278780
rect 329064 278740 329070 278752
rect 329190 278740 329196 278752
rect 329248 278740 329254 278792
rect 335814 278740 335820 278792
rect 335872 278780 335878 278792
rect 335998 278780 336004 278792
rect 335872 278752 336004 278780
rect 335872 278740 335878 278752
rect 335998 278740 336004 278752
rect 336056 278740 336062 278792
rect 264514 278712 264520 278724
rect 264475 278684 264520 278712
rect 264514 278672 264520 278684
rect 264572 278672 264578 278724
rect 265802 278712 265808 278724
rect 265763 278684 265808 278712
rect 265802 278672 265808 278684
rect 265860 278672 265866 278724
rect 258718 277420 258724 277432
rect 258679 277392 258724 277420
rect 258718 277380 258724 277392
rect 258776 277380 258782 277432
rect 232682 273300 232688 273352
rect 232740 273300 232746 273352
rect 341610 273300 341616 273352
rect 341668 273300 341674 273352
rect 232700 273216 232728 273300
rect 260282 273272 260288 273284
rect 260243 273244 260288 273272
rect 260282 273232 260288 273244
rect 260340 273232 260346 273284
rect 333146 273272 333152 273284
rect 333072 273244 333152 273272
rect 333072 273216 333100 273244
rect 333146 273232 333152 273244
rect 333204 273232 333210 273284
rect 341628 273216 341656 273300
rect 232682 273164 232688 273216
rect 232740 273164 232746 273216
rect 333054 273164 333060 273216
rect 333112 273164 333118 273216
rect 341610 273164 341616 273216
rect 341668 273164 341674 273216
rect 246482 272552 246488 272604
rect 246540 272592 246546 272604
rect 246758 272592 246764 272604
rect 246540 272564 246764 272592
rect 246540 272552 246546 272564
rect 246758 272552 246764 272564
rect 246816 272552 246822 272604
rect 328914 270580 328920 270632
rect 328972 270580 328978 270632
rect 231210 270552 231216 270564
rect 231171 270524 231216 270552
rect 231210 270512 231216 270524
rect 231268 270512 231274 270564
rect 240686 270552 240692 270564
rect 240647 270524 240692 270552
rect 240686 270512 240692 270524
rect 240744 270512 240750 270564
rect 246022 270552 246028 270564
rect 245983 270524 246028 270552
rect 246022 270512 246028 270524
rect 246080 270512 246086 270564
rect 328932 270496 328960 270580
rect 345290 270512 345296 270564
rect 345348 270552 345354 270564
rect 345382 270552 345388 270564
rect 345348 270524 345388 270552
rect 345348 270512 345354 270524
rect 345382 270512 345388 270524
rect 345440 270512 345446 270564
rect 100662 270484 100668 270496
rect 100623 270456 100668 270484
rect 100662 270444 100668 270456
rect 100720 270444 100726 270496
rect 238018 270484 238024 270496
rect 237979 270456 238024 270484
rect 238018 270444 238024 270456
rect 238076 270444 238082 270496
rect 244918 270444 244924 270496
rect 244976 270484 244982 270496
rect 245102 270484 245108 270496
rect 244976 270456 245108 270484
rect 244976 270444 244982 270456
rect 245102 270444 245108 270456
rect 245160 270444 245166 270496
rect 328914 270444 328920 270496
rect 328972 270444 328978 270496
rect 107470 269084 107476 269136
rect 107528 269124 107534 269136
rect 107654 269124 107660 269136
rect 107528 269096 107660 269124
rect 107528 269084 107534 269096
rect 107654 269084 107660 269096
rect 107712 269084 107718 269136
rect 231946 269084 231952 269136
rect 232004 269124 232010 269136
rect 232130 269124 232136 269136
rect 232004 269096 232136 269124
rect 232004 269084 232010 269096
rect 232130 269084 232136 269096
rect 232188 269084 232194 269136
rect 261386 269084 261392 269136
rect 261444 269124 261450 269136
rect 261662 269124 261668 269136
rect 261444 269096 261668 269124
rect 261444 269084 261450 269096
rect 261662 269084 261668 269096
rect 261720 269084 261726 269136
rect 264514 269124 264520 269136
rect 264475 269096 264520 269124
rect 264514 269084 264520 269096
rect 264572 269084 264578 269136
rect 265802 269124 265808 269136
rect 265763 269096 265808 269124
rect 265802 269084 265808 269096
rect 265860 269084 265866 269136
rect 320910 269084 320916 269136
rect 320968 269124 320974 269136
rect 321094 269124 321100 269136
rect 320968 269096 321100 269124
rect 320968 269084 320974 269096
rect 321094 269084 321100 269096
rect 321152 269084 321158 269136
rect 319438 267724 319444 267776
rect 319496 267764 319502 267776
rect 319622 267764 319628 267776
rect 319496 267736 319628 267764
rect 319496 267724 319502 267736
rect 319622 267724 319628 267736
rect 319680 267724 319686 267776
rect 326338 267724 326344 267776
rect 326396 267764 326402 267776
rect 326522 267764 326528 267776
rect 326396 267736 326528 267764
rect 326396 267724 326402 267736
rect 326522 267724 326528 267736
rect 326580 267724 326586 267776
rect 331582 266296 331588 266348
rect 331640 266336 331646 266348
rect 331858 266336 331864 266348
rect 331640 266308 331864 266336
rect 331640 266296 331646 266308
rect 331858 266296 331864 266308
rect 331916 266296 331922 266348
rect 2774 266092 2780 266144
rect 2832 266132 2838 266144
rect 5350 266132 5356 266144
rect 2832 266104 5356 266132
rect 2832 266092 2838 266104
rect 5350 266092 5356 266104
rect 5408 266092 5414 266144
rect 260285 265319 260343 265325
rect 260285 265285 260297 265319
rect 260331 265316 260343 265319
rect 260374 265316 260380 265328
rect 260331 265288 260380 265316
rect 260331 265285 260343 265288
rect 260285 265279 260343 265285
rect 260374 265276 260380 265288
rect 260432 265276 260438 265328
rect 322290 263616 322296 263628
rect 322251 263588 322296 263616
rect 322290 263576 322296 263588
rect 322348 263576 322354 263628
rect 333054 263576 333060 263628
rect 333112 263576 333118 263628
rect 333072 263548 333100 263576
rect 333146 263548 333152 263560
rect 333072 263520 333152 263548
rect 333146 263508 333152 263520
rect 333204 263508 333210 263560
rect 231762 262896 231768 262948
rect 231820 262936 231826 262948
rect 232038 262936 232044 262948
rect 231820 262908 232044 262936
rect 231820 262896 231826 262908
rect 232038 262896 232044 262908
rect 232096 262896 232102 262948
rect 100662 260896 100668 260908
rect 100623 260868 100668 260896
rect 100662 260856 100668 260868
rect 100720 260856 100726 260908
rect 238018 260896 238024 260908
rect 237979 260868 238024 260896
rect 238018 260856 238024 260868
rect 238076 260856 238082 260908
rect 328914 260856 328920 260908
rect 328972 260896 328978 260908
rect 329006 260896 329012 260908
rect 328972 260868 329012 260896
rect 328972 260856 328978 260868
rect 329006 260856 329012 260868
rect 329064 260856 329070 260908
rect 333238 260856 333244 260908
rect 333296 260896 333302 260908
rect 333330 260896 333336 260908
rect 333296 260868 333336 260896
rect 333296 260856 333302 260868
rect 333330 260856 333336 260868
rect 333388 260856 333394 260908
rect 334526 260856 334532 260908
rect 334584 260896 334590 260908
rect 334618 260896 334624 260908
rect 334584 260868 334624 260896
rect 334584 260856 334590 260868
rect 334618 260856 334624 260868
rect 334676 260856 334682 260908
rect 335722 260856 335728 260908
rect 335780 260896 335786 260908
rect 335814 260896 335820 260908
rect 335780 260868 335820 260896
rect 335780 260856 335786 260868
rect 335814 260856 335820 260868
rect 335872 260856 335878 260908
rect 231210 260828 231216 260840
rect 231171 260800 231216 260828
rect 231210 260788 231216 260800
rect 231268 260788 231274 260840
rect 330478 260788 330484 260840
rect 330536 260828 330542 260840
rect 330570 260828 330576 260840
rect 330536 260800 330576 260828
rect 330536 260788 330542 260800
rect 330570 260788 330576 260800
rect 330628 260788 330634 260840
rect 341610 260828 341616 260840
rect 341571 260800 341616 260828
rect 341610 260788 341616 260800
rect 341668 260788 341674 260840
rect 345382 260788 345388 260840
rect 345440 260788 345446 260840
rect 345400 260704 345428 260788
rect 345382 260652 345388 260704
rect 345440 260652 345446 260704
rect 257062 259428 257068 259480
rect 257120 259468 257126 259480
rect 257154 259468 257160 259480
rect 257120 259440 257160 259468
rect 257120 259428 257126 259440
rect 257154 259428 257160 259440
rect 257212 259428 257218 259480
rect 264330 259428 264336 259480
rect 264388 259468 264394 259480
rect 264514 259468 264520 259480
rect 264388 259440 264520 259468
rect 264388 259428 264394 259440
rect 264514 259428 264520 259440
rect 264572 259428 264578 259480
rect 265618 259428 265624 259480
rect 265676 259468 265682 259480
rect 265802 259468 265808 259480
rect 265676 259440 265808 259468
rect 265676 259428 265682 259440
rect 265802 259428 265808 259440
rect 265860 259428 265866 259480
rect 293126 259428 293132 259480
rect 293184 259468 293190 259480
rect 293310 259468 293316 259480
rect 293184 259440 293316 259468
rect 293184 259428 293190 259440
rect 293310 259428 293316 259440
rect 293368 259428 293374 259480
rect 320910 259428 320916 259480
rect 320968 259468 320974 259480
rect 321094 259468 321100 259480
rect 320968 259440 321100 259468
rect 320968 259428 320974 259440
rect 321094 259428 321100 259440
rect 321152 259428 321158 259480
rect 322290 259468 322296 259480
rect 322251 259440 322296 259468
rect 322290 259428 322296 259440
rect 322348 259428 322354 259480
rect 244918 259360 244924 259412
rect 244976 259400 244982 259412
rect 245102 259400 245108 259412
rect 244976 259372 245108 259400
rect 244976 259360 244982 259372
rect 245102 259360 245108 259372
rect 245160 259360 245166 259412
rect 246298 258068 246304 258120
rect 246356 258108 246362 258120
rect 246390 258108 246396 258120
rect 246356 258080 246396 258108
rect 246356 258068 246362 258080
rect 246390 258068 246396 258080
rect 246448 258068 246454 258120
rect 258626 258068 258632 258120
rect 258684 258108 258690 258120
rect 258718 258108 258724 258120
rect 258684 258080 258724 258108
rect 258684 258068 258690 258080
rect 258718 258068 258724 258080
rect 258776 258068 258782 258120
rect 232038 258000 232044 258052
rect 232096 258040 232102 258052
rect 232133 258043 232191 258049
rect 232133 258040 232145 258043
rect 232096 258012 232145 258040
rect 232096 258000 232102 258012
rect 232133 258009 232145 258012
rect 232179 258009 232191 258043
rect 232133 258003 232191 258009
rect 232314 258000 232320 258052
rect 232372 258040 232378 258052
rect 232409 258043 232467 258049
rect 232409 258040 232421 258043
rect 232372 258012 232421 258040
rect 232372 258000 232378 258012
rect 232409 258009 232421 258012
rect 232455 258009 232467 258043
rect 244366 258040 244372 258052
rect 244327 258012 244372 258040
rect 232409 258003 232467 258009
rect 244366 258000 244372 258012
rect 244424 258000 244430 258052
rect 319622 258040 319628 258052
rect 319583 258012 319628 258040
rect 319622 258000 319628 258012
rect 319680 258000 319686 258052
rect 322106 258000 322112 258052
rect 322164 258040 322170 258052
rect 322198 258040 322204 258052
rect 322164 258012 322204 258040
rect 322164 258000 322170 258012
rect 322198 258000 322204 258012
rect 322256 258000 322262 258052
rect 335725 258043 335783 258049
rect 335725 258009 335737 258043
rect 335771 258040 335783 258043
rect 335814 258040 335820 258052
rect 335771 258012 335820 258040
rect 335771 258009 335783 258012
rect 335725 258003 335783 258009
rect 335814 258000 335820 258012
rect 335872 258000 335878 258052
rect 299014 256680 299020 256692
rect 298975 256652 299020 256680
rect 299014 256640 299020 256652
rect 299072 256640 299078 256692
rect 334526 256680 334532 256692
rect 334487 256652 334532 256680
rect 334526 256640 334532 256652
rect 334584 256640 334590 256692
rect 326249 254099 326307 254105
rect 326249 254065 326261 254099
rect 326295 254096 326307 254099
rect 326338 254096 326344 254108
rect 326295 254068 326344 254096
rect 326295 254065 326307 254068
rect 326249 254059 326307 254065
rect 326338 254056 326344 254068
rect 326396 254056 326402 254108
rect 253106 254028 253112 254040
rect 253032 254000 253112 254028
rect 253032 253904 253060 254000
rect 253106 253988 253112 254000
rect 253164 253988 253170 254040
rect 333146 253960 333152 253972
rect 333072 253932 333152 253960
rect 333072 253904 333100 253932
rect 333146 253920 333152 253932
rect 333204 253920 333210 253972
rect 232130 253892 232136 253904
rect 232091 253864 232136 253892
rect 232130 253852 232136 253864
rect 232188 253852 232194 253904
rect 253014 253852 253020 253904
rect 253072 253852 253078 253904
rect 333054 253852 333060 253904
rect 333112 253852 333118 253904
rect 232314 253172 232320 253224
rect 232372 253212 232378 253224
rect 232409 253215 232467 253221
rect 232409 253212 232421 253215
rect 232372 253184 232421 253212
rect 232372 253172 232378 253184
rect 232409 253181 232421 253184
rect 232455 253181 232467 253215
rect 232409 253175 232467 253181
rect 265618 253172 265624 253224
rect 265676 253212 265682 253224
rect 265802 253212 265808 253224
rect 265676 253184 265808 253212
rect 265676 253172 265682 253184
rect 265802 253172 265808 253184
rect 265860 253172 265866 253224
rect 231210 251240 231216 251252
rect 231171 251212 231216 251240
rect 231210 251200 231216 251212
rect 231268 251200 231274 251252
rect 256970 251240 256976 251252
rect 256931 251212 256976 251240
rect 256970 251200 256976 251212
rect 257028 251200 257034 251252
rect 341613 251243 341671 251249
rect 341613 251209 341625 251243
rect 341659 251240 341671 251243
rect 341702 251240 341708 251252
rect 341659 251212 341708 251240
rect 341659 251209 341671 251212
rect 341613 251203 341671 251209
rect 341702 251200 341708 251212
rect 341760 251200 341766 251252
rect 100662 251172 100668 251184
rect 100623 251144 100668 251172
rect 100662 251132 100668 251144
rect 100720 251132 100726 251184
rect 334526 251104 334532 251116
rect 334487 251076 334532 251104
rect 334526 251064 334532 251076
rect 334584 251064 334590 251116
rect 335725 250971 335783 250977
rect 335725 250937 335737 250971
rect 335771 250968 335783 250971
rect 335814 250968 335820 250980
rect 335771 250940 335820 250968
rect 335771 250937 335783 250940
rect 335725 250931 335783 250937
rect 335814 250928 335820 250940
rect 335872 250928 335878 250980
rect 258626 249840 258632 249892
rect 258684 249840 258690 249892
rect 107470 249772 107476 249824
rect 107528 249812 107534 249824
rect 107654 249812 107660 249824
rect 107528 249784 107660 249812
rect 107528 249772 107534 249784
rect 107654 249772 107660 249784
rect 107712 249772 107718 249824
rect 256970 249812 256976 249824
rect 256931 249784 256976 249812
rect 256970 249772 256976 249784
rect 257028 249772 257034 249824
rect 258644 249812 258672 249840
rect 258718 249812 258724 249824
rect 258644 249784 258724 249812
rect 258718 249772 258724 249784
rect 258776 249772 258782 249824
rect 320910 249772 320916 249824
rect 320968 249812 320974 249824
rect 321094 249812 321100 249824
rect 320968 249784 321100 249812
rect 320968 249772 320974 249784
rect 321094 249772 321100 249784
rect 321152 249772 321158 249824
rect 326246 249812 326252 249824
rect 326207 249784 326252 249812
rect 326246 249772 326252 249784
rect 326304 249772 326310 249824
rect 345382 249772 345388 249824
rect 345440 249812 345446 249824
rect 345566 249812 345572 249824
rect 345440 249784 345572 249812
rect 345440 249772 345446 249784
rect 345566 249772 345572 249784
rect 345624 249772 345630 249824
rect 258810 249744 258816 249756
rect 258771 249716 258816 249744
rect 258810 249704 258816 249716
rect 258868 249704 258874 249756
rect 246298 248384 246304 248396
rect 246259 248356 246304 248384
rect 246298 248344 246304 248356
rect 246356 248344 246362 248396
rect 299014 247092 299020 247104
rect 298975 247064 299020 247092
rect 299014 247052 299020 247064
rect 299072 247052 299078 247104
rect 300302 247024 300308 247036
rect 300263 246996 300308 247024
rect 300302 246984 300308 246996
rect 300360 246984 300366 247036
rect 301774 247024 301780 247036
rect 301735 246996 301780 247024
rect 301774 246984 301780 246996
rect 301832 246984 301838 247036
rect 330478 246984 330484 247036
rect 330536 247024 330542 247036
rect 330570 247024 330576 247036
rect 330536 246996 330576 247024
rect 330536 246984 330542 246996
rect 330570 246984 330576 246996
rect 330628 246984 330634 247036
rect 331766 246984 331772 247036
rect 331824 247024 331830 247036
rect 331950 247024 331956 247036
rect 331824 246996 331956 247024
rect 331824 246984 331830 246996
rect 331950 246984 331956 246996
rect 332008 246984 332014 247036
rect 333238 246984 333244 247036
rect 333296 247024 333302 247036
rect 333422 247024 333428 247036
rect 333296 246996 333428 247024
rect 333296 246984 333302 246996
rect 333422 246984 333428 246996
rect 333480 246984 333486 247036
rect 333054 244264 333060 244316
rect 333112 244264 333118 244316
rect 340046 244264 340052 244316
rect 340104 244264 340110 244316
rect 344094 244264 344100 244316
rect 344152 244304 344158 244316
rect 344278 244304 344284 244316
rect 344152 244276 344284 244304
rect 344152 244264 344158 244276
rect 344278 244264 344284 244276
rect 344336 244264 344342 244316
rect 333072 244236 333100 244264
rect 333146 244236 333152 244248
rect 333072 244208 333152 244236
rect 333146 244196 333152 244208
rect 333204 244196 333210 244248
rect 340064 244168 340092 244264
rect 340138 244168 340144 244180
rect 340064 244140 340144 244168
rect 340138 244128 340144 244140
rect 340196 244128 340202 244180
rect 244366 241584 244372 241596
rect 244327 241556 244372 241584
rect 244366 241544 244372 241556
rect 244424 241544 244430 241596
rect 100662 241516 100668 241528
rect 100623 241488 100668 241516
rect 100662 241476 100668 241488
rect 100720 241476 100726 241528
rect 253014 241476 253020 241528
rect 253072 241516 253078 241528
rect 253106 241516 253112 241528
rect 253072 241488 253112 241516
rect 253072 241476 253078 241488
rect 253106 241476 253112 241488
rect 253164 241476 253170 241528
rect 335814 241476 335820 241528
rect 335872 241516 335878 241528
rect 335998 241516 336004 241528
rect 335872 241488 336004 241516
rect 335872 241476 335878 241488
rect 335998 241476 336004 241488
rect 336056 241476 336062 241528
rect 260190 240252 260196 240304
rect 260248 240292 260254 240304
rect 260248 240264 260328 240292
rect 260248 240252 260254 240264
rect 258810 240224 258816 240236
rect 258771 240196 258816 240224
rect 258810 240184 258816 240196
rect 258868 240184 258874 240236
rect 260300 240168 260328 240264
rect 232038 240116 232044 240168
rect 232096 240156 232102 240168
rect 232130 240156 232136 240168
rect 232096 240128 232136 240156
rect 232096 240116 232102 240128
rect 232130 240116 232136 240128
rect 232188 240116 232194 240168
rect 260282 240116 260288 240168
rect 260340 240116 260346 240168
rect 261478 240116 261484 240168
rect 261536 240156 261542 240168
rect 261570 240156 261576 240168
rect 261536 240128 261576 240156
rect 261536 240116 261542 240128
rect 261570 240116 261576 240128
rect 261628 240116 261634 240168
rect 264330 240116 264336 240168
rect 264388 240156 264394 240168
rect 264514 240156 264520 240168
rect 264388 240128 264520 240156
rect 264388 240116 264394 240128
rect 264514 240116 264520 240128
rect 264572 240116 264578 240168
rect 293126 240116 293132 240168
rect 293184 240156 293190 240168
rect 293310 240156 293316 240168
rect 293184 240128 293316 240156
rect 293184 240116 293190 240128
rect 293310 240116 293316 240128
rect 293368 240116 293374 240168
rect 319622 240156 319628 240168
rect 319583 240128 319628 240156
rect 319622 240116 319628 240128
rect 319680 240116 319686 240168
rect 320910 240116 320916 240168
rect 320968 240156 320974 240168
rect 321094 240156 321100 240168
rect 320968 240128 321100 240156
rect 320968 240116 320974 240128
rect 321094 240116 321100 240128
rect 321152 240116 321158 240168
rect 232682 240088 232688 240100
rect 232643 240060 232688 240088
rect 232682 240048 232688 240060
rect 232740 240048 232746 240100
rect 258626 240048 258632 240100
rect 258684 240088 258690 240100
rect 258810 240088 258816 240100
rect 258684 240060 258816 240088
rect 258684 240048 258690 240060
rect 258810 240048 258816 240060
rect 258868 240048 258874 240100
rect 246301 238799 246359 238805
rect 246301 238765 246313 238799
rect 246347 238796 246359 238799
rect 246390 238796 246396 238808
rect 246347 238768 246396 238796
rect 246347 238765 246359 238768
rect 246301 238759 246359 238765
rect 246390 238756 246396 238768
rect 246448 238756 246454 238808
rect 261570 238728 261576 238740
rect 261531 238700 261576 238728
rect 261570 238688 261576 238700
rect 261628 238688 261634 238740
rect 265618 238688 265624 238740
rect 265676 238728 265682 238740
rect 265802 238728 265808 238740
rect 265676 238700 265808 238728
rect 265676 238688 265682 238700
rect 265802 238688 265808 238700
rect 265860 238688 265866 238740
rect 319438 238688 319444 238740
rect 319496 238728 319502 238740
rect 319622 238728 319628 238740
rect 319496 238700 319628 238728
rect 319496 238688 319502 238700
rect 319622 238688 319628 238700
rect 319680 238688 319686 238740
rect 322106 238688 322112 238740
rect 322164 238728 322170 238740
rect 322290 238728 322296 238740
rect 322164 238700 322296 238728
rect 322164 238688 322170 238700
rect 322290 238688 322296 238700
rect 322348 238688 322354 238740
rect 300302 237436 300308 237448
rect 300263 237408 300308 237436
rect 300302 237396 300308 237408
rect 300360 237396 300366 237448
rect 301774 237436 301780 237448
rect 301735 237408 301780 237436
rect 301774 237396 301780 237408
rect 301832 237396 301838 237448
rect 299014 237368 299020 237380
rect 298975 237340 299020 237368
rect 299014 237328 299020 237340
rect 299072 237328 299078 237380
rect 329006 237328 329012 237380
rect 329064 237368 329070 237380
rect 329190 237368 329196 237380
rect 329064 237340 329196 237368
rect 329064 237328 329070 237340
rect 329190 237328 329196 237340
rect 329248 237328 329254 237380
rect 330386 237328 330392 237380
rect 330444 237368 330450 237380
rect 330478 237368 330484 237380
rect 330444 237340 330484 237368
rect 330444 237328 330450 237340
rect 330478 237328 330484 237340
rect 330536 237328 330542 237380
rect 2774 237260 2780 237312
rect 2832 237300 2838 237312
rect 5258 237300 5264 237312
rect 2832 237272 5264 237300
rect 2832 237260 2838 237272
rect 5258 237260 5264 237272
rect 5316 237260 5322 237312
rect 301774 235940 301780 235952
rect 301735 235912 301780 235940
rect 301774 235900 301780 235912
rect 301832 235900 301838 235952
rect 330386 235940 330392 235952
rect 330347 235912 330392 235940
rect 330386 235900 330392 235912
rect 330444 235900 330450 235952
rect 232682 235328 232688 235340
rect 232643 235300 232688 235328
rect 232682 235288 232688 235300
rect 232740 235288 232746 235340
rect 232038 234648 232044 234660
rect 231999 234620 232044 234648
rect 232038 234608 232044 234620
rect 232096 234608 232102 234660
rect 245010 234648 245016 234660
rect 244936 234620 245016 234648
rect 244936 234592 244964 234620
rect 245010 234608 245016 234620
rect 245068 234608 245074 234660
rect 246390 234608 246396 234660
rect 246448 234608 246454 234660
rect 244182 234540 244188 234592
rect 244240 234580 244246 234592
rect 244366 234580 244372 234592
rect 244240 234552 244372 234580
rect 244240 234540 244246 234552
rect 244366 234540 244372 234552
rect 244424 234540 244430 234592
rect 244918 234540 244924 234592
rect 244976 234540 244982 234592
rect 246408 234512 246436 234608
rect 261570 234580 261576 234592
rect 261531 234552 261576 234580
rect 261570 234540 261576 234552
rect 261628 234540 261634 234592
rect 246482 234512 246488 234524
rect 246408 234484 246488 234512
rect 246482 234472 246488 234484
rect 246540 234472 246546 234524
rect 231210 231820 231216 231872
rect 231268 231860 231274 231872
rect 231394 231860 231400 231872
rect 231268 231832 231400 231860
rect 231268 231820 231274 231832
rect 231394 231820 231400 231832
rect 231452 231820 231458 231872
rect 331766 231820 331772 231872
rect 331824 231820 331830 231872
rect 335814 231820 335820 231872
rect 335872 231820 335878 231872
rect 331784 231792 331812 231820
rect 331858 231792 331864 231804
rect 331784 231764 331864 231792
rect 331858 231752 331864 231764
rect 331916 231752 331922 231804
rect 335832 231792 335860 231820
rect 335906 231792 335912 231804
rect 335832 231764 335912 231792
rect 335906 231752 335912 231764
rect 335964 231752 335970 231804
rect 253014 230528 253020 230580
rect 253072 230568 253078 230580
rect 253106 230568 253112 230580
rect 253072 230540 253112 230568
rect 253072 230528 253078 230540
rect 253106 230528 253112 230540
rect 253164 230528 253170 230580
rect 340138 230528 340144 230580
rect 340196 230528 340202 230580
rect 107470 230460 107476 230512
rect 107528 230500 107534 230512
rect 107654 230500 107660 230512
rect 107528 230472 107660 230500
rect 107528 230460 107534 230472
rect 107654 230460 107660 230472
rect 107712 230460 107718 230512
rect 232038 230500 232044 230512
rect 231999 230472 232044 230500
rect 232038 230460 232044 230472
rect 232096 230460 232102 230512
rect 237834 230460 237840 230512
rect 237892 230500 237898 230512
rect 237926 230500 237932 230512
rect 237892 230472 237932 230500
rect 237892 230460 237898 230472
rect 237926 230460 237932 230472
rect 237984 230460 237990 230512
rect 240502 230460 240508 230512
rect 240560 230500 240566 230512
rect 240686 230500 240692 230512
rect 240560 230472 240692 230500
rect 240560 230460 240566 230472
rect 240686 230460 240692 230472
rect 240744 230460 240750 230512
rect 257062 230460 257068 230512
rect 257120 230500 257126 230512
rect 257154 230500 257160 230512
rect 257120 230472 257160 230500
rect 257120 230460 257126 230472
rect 257154 230460 257160 230472
rect 257212 230460 257218 230512
rect 320910 230460 320916 230512
rect 320968 230500 320974 230512
rect 321094 230500 321100 230512
rect 320968 230472 321100 230500
rect 320968 230460 320974 230472
rect 321094 230460 321100 230472
rect 321152 230460 321158 230512
rect 326246 230460 326252 230512
rect 326304 230500 326310 230512
rect 326338 230500 326344 230512
rect 326304 230472 326344 230500
rect 326304 230460 326310 230472
rect 326338 230460 326344 230472
rect 326396 230460 326402 230512
rect 339954 230460 339960 230512
rect 340012 230500 340018 230512
rect 340156 230500 340184 230528
rect 340012 230472 340184 230500
rect 340012 230460 340018 230472
rect 330389 230095 330447 230101
rect 330389 230061 330401 230095
rect 330435 230092 330447 230095
rect 330754 230092 330760 230104
rect 330435 230064 330760 230092
rect 330435 230061 330447 230064
rect 330389 230055 330447 230061
rect 330754 230052 330760 230064
rect 330812 230052 330818 230104
rect 260190 229168 260196 229220
rect 260248 229208 260254 229220
rect 260374 229208 260380 229220
rect 260248 229180 260380 229208
rect 260248 229168 260254 229180
rect 260374 229168 260380 229180
rect 260432 229168 260438 229220
rect 260374 229072 260380 229084
rect 260335 229044 260380 229072
rect 260374 229032 260380 229044
rect 260432 229032 260438 229084
rect 340049 229075 340107 229081
rect 340049 229041 340061 229075
rect 340095 229072 340107 229075
rect 340138 229072 340144 229084
rect 340095 229044 340144 229072
rect 340095 229041 340107 229044
rect 340049 229035 340107 229041
rect 340138 229032 340144 229044
rect 340196 229032 340202 229084
rect 299014 227780 299020 227792
rect 298975 227752 299020 227780
rect 299014 227740 299020 227752
rect 299072 227740 299078 227792
rect 300302 227712 300308 227724
rect 300263 227684 300308 227712
rect 300302 227672 300308 227684
rect 300360 227672 300366 227724
rect 333054 227712 333060 227724
rect 333015 227684 333060 227712
rect 333054 227672 333060 227684
rect 333112 227672 333118 227724
rect 299014 227644 299020 227656
rect 298975 227616 299020 227644
rect 299014 227604 299020 227616
rect 299072 227604 299078 227656
rect 267182 227060 267188 227112
rect 267240 227060 267246 227112
rect 268654 227060 268660 227112
rect 268712 227060 268718 227112
rect 267200 226976 267228 227060
rect 268672 226976 268700 227060
rect 267182 226924 267188 226976
rect 267240 226924 267246 226976
rect 268654 226924 268660 226976
rect 268712 226924 268718 226976
rect 301774 226352 301780 226364
rect 301735 226324 301780 226352
rect 301774 226312 301780 226324
rect 301832 226312 301838 226364
rect 232038 224992 232044 225004
rect 231999 224964 232044 224992
rect 232038 224952 232044 224964
rect 232096 224952 232102 225004
rect 257062 224952 257068 225004
rect 257120 224992 257126 225004
rect 257120 224964 257200 224992
rect 257120 224952 257126 224964
rect 257172 224936 257200 224964
rect 344094 224952 344100 225004
rect 344152 224992 344158 225004
rect 344278 224992 344284 225004
rect 344152 224964 344284 224992
rect 344152 224952 344158 224964
rect 344278 224952 344284 224964
rect 344336 224952 344342 225004
rect 257154 224884 257160 224936
rect 257212 224884 257218 224936
rect 330754 224884 330760 224936
rect 330812 224924 330818 224936
rect 330938 224924 330944 224936
rect 330812 224896 330944 224924
rect 330812 224884 330818 224896
rect 330938 224884 330944 224896
rect 330996 224884 331002 224936
rect 260374 224244 260380 224256
rect 260335 224216 260380 224244
rect 260374 224204 260380 224216
rect 260432 224204 260438 224256
rect 322106 224204 322112 224256
rect 322164 224244 322170 224256
rect 322290 224244 322296 224256
rect 322164 224216 322296 224244
rect 322164 224204 322170 224216
rect 322290 224204 322296 224216
rect 322348 224204 322354 224256
rect 2774 223048 2780 223100
rect 2832 223088 2838 223100
rect 5166 223088 5172 223100
rect 2832 223060 5172 223088
rect 2832 223048 2838 223060
rect 5166 223048 5172 223060
rect 5224 223048 5230 223100
rect 232314 222232 232320 222284
rect 232372 222272 232378 222284
rect 232590 222272 232596 222284
rect 232372 222244 232596 222272
rect 232372 222232 232378 222244
rect 232590 222232 232596 222244
rect 232648 222232 232654 222284
rect 100662 222164 100668 222216
rect 100720 222204 100726 222216
rect 100846 222204 100852 222216
rect 100720 222176 100852 222204
rect 100720 222164 100726 222176
rect 100846 222164 100852 222176
rect 100904 222164 100910 222216
rect 232038 222204 232044 222216
rect 231999 222176 232044 222204
rect 232038 222164 232044 222176
rect 232096 222164 232102 222216
rect 237926 222164 237932 222216
rect 237984 222204 237990 222216
rect 238018 222204 238024 222216
rect 237984 222176 238024 222204
rect 237984 222164 237990 222176
rect 238018 222164 238024 222176
rect 238076 222164 238082 222216
rect 331766 222164 331772 222216
rect 331824 222204 331830 222216
rect 331858 222204 331864 222216
rect 331824 222176 331864 222204
rect 331824 222164 331830 222176
rect 331858 222164 331864 222176
rect 331916 222164 331922 222216
rect 333238 222164 333244 222216
rect 333296 222204 333302 222216
rect 333330 222204 333336 222216
rect 333296 222176 333336 222204
rect 333296 222164 333302 222176
rect 333330 222164 333336 222176
rect 333388 222164 333394 222216
rect 326338 220912 326344 220924
rect 326264 220884 326344 220912
rect 326264 220856 326292 220884
rect 326338 220872 326344 220884
rect 326396 220872 326402 220924
rect 253106 220804 253112 220856
rect 253164 220844 253170 220856
rect 253290 220844 253296 220856
rect 253164 220816 253296 220844
rect 253164 220804 253170 220816
rect 253290 220804 253296 220816
rect 253348 220804 253354 220856
rect 293126 220804 293132 220856
rect 293184 220844 293190 220856
rect 293310 220844 293316 220856
rect 293184 220816 293316 220844
rect 293184 220804 293190 220816
rect 293310 220804 293316 220816
rect 293368 220804 293374 220856
rect 320910 220804 320916 220856
rect 320968 220844 320974 220856
rect 321094 220844 321100 220856
rect 320968 220816 321100 220844
rect 320968 220804 320974 220816
rect 321094 220804 321100 220816
rect 321152 220804 321158 220856
rect 326246 220804 326252 220856
rect 326304 220804 326310 220856
rect 340046 220776 340052 220788
rect 340007 220748 340052 220776
rect 340046 220736 340052 220748
rect 340104 220736 340110 220788
rect 260374 219416 260380 219428
rect 260335 219388 260380 219416
rect 260374 219376 260380 219388
rect 260432 219376 260438 219428
rect 261570 219416 261576 219428
rect 261531 219388 261576 219416
rect 261570 219376 261576 219388
rect 261628 219376 261634 219428
rect 265618 219376 265624 219428
rect 265676 219416 265682 219428
rect 265802 219416 265808 219428
rect 265676 219388 265808 219416
rect 265676 219376 265682 219388
rect 265802 219376 265808 219388
rect 265860 219376 265866 219428
rect 319622 219416 319628 219428
rect 319583 219388 319628 219416
rect 319622 219376 319628 219388
rect 319680 219376 319686 219428
rect 321094 219416 321100 219428
rect 321055 219388 321100 219416
rect 321094 219376 321100 219388
rect 321152 219376 321158 219428
rect 322109 219351 322167 219357
rect 322109 219317 322121 219351
rect 322155 219348 322167 219351
rect 322290 219348 322296 219360
rect 322155 219320 322296 219348
rect 322155 219317 322167 219320
rect 322109 219311 322167 219317
rect 322290 219308 322296 219320
rect 322348 219308 322354 219360
rect 299014 218056 299020 218068
rect 298975 218028 299020 218056
rect 299014 218016 299020 218028
rect 299072 218016 299078 218068
rect 300302 218056 300308 218068
rect 300263 218028 300308 218056
rect 300302 218016 300308 218028
rect 300360 218016 300366 218068
rect 333057 218059 333115 218065
rect 333057 218025 333069 218059
rect 333103 218056 333115 218059
rect 333146 218056 333152 218068
rect 333103 218028 333152 218056
rect 333103 218025 333115 218028
rect 333057 218019 333115 218025
rect 333146 218016 333152 218028
rect 333204 218016 333210 218068
rect 335814 218016 335820 218068
rect 335872 218056 335878 218068
rect 335906 218056 335912 218068
rect 335872 218028 335912 218056
rect 335872 218016 335878 218028
rect 335906 218016 335912 218028
rect 335964 218016 335970 218068
rect 333238 217948 333244 218000
rect 333296 217948 333302 218000
rect 333256 217920 333284 217948
rect 333330 217920 333336 217932
rect 333256 217892 333336 217920
rect 333330 217880 333336 217892
rect 333388 217880 333394 217932
rect 246393 217447 246451 217453
rect 246393 217413 246405 217447
rect 246439 217444 246451 217447
rect 246482 217444 246488 217456
rect 246439 217416 246488 217444
rect 246439 217413 246451 217416
rect 246393 217407 246451 217413
rect 246482 217404 246488 217416
rect 246540 217404 246546 217456
rect 301774 216628 301780 216640
rect 301735 216600 301780 216628
rect 301774 216588 301780 216600
rect 301832 216588 301838 216640
rect 334526 216588 334532 216640
rect 334584 216628 334590 216640
rect 334621 216631 334679 216637
rect 334621 216628 334633 216631
rect 334584 216600 334633 216628
rect 334584 216588 334590 216600
rect 334621 216597 334633 216600
rect 334667 216597 334679 216631
rect 334621 216591 334679 216597
rect 341702 215976 341708 216028
rect 341760 216016 341766 216028
rect 341886 216016 341892 216028
rect 341760 215988 341892 216016
rect 341760 215976 341766 215988
rect 341886 215976 341892 215988
rect 341944 215976 341950 216028
rect 326246 215404 326252 215416
rect 326207 215376 326252 215404
rect 326246 215364 326252 215376
rect 326304 215364 326310 215416
rect 261570 215268 261576 215280
rect 261531 215240 261576 215268
rect 261570 215228 261576 215240
rect 261628 215228 261634 215280
rect 329006 215268 329012 215280
rect 328967 215240 329012 215268
rect 329006 215228 329012 215240
rect 329064 215228 329070 215280
rect 330754 215228 330760 215280
rect 330812 215268 330818 215280
rect 330938 215268 330944 215280
rect 330812 215240 330944 215268
rect 330812 215228 330818 215240
rect 330938 215228 330944 215240
rect 330996 215228 331002 215280
rect 232590 215092 232596 215144
rect 232648 215132 232654 215144
rect 232774 215132 232780 215144
rect 232648 215104 232780 215132
rect 232648 215092 232654 215104
rect 232774 215092 232780 215104
rect 232832 215092 232838 215144
rect 260374 214520 260380 214532
rect 260335 214492 260380 214520
rect 260374 214480 260380 214492
rect 260432 214480 260438 214532
rect 245010 212644 245016 212696
rect 245068 212644 245074 212696
rect 231210 212508 231216 212560
rect 231268 212548 231274 212560
rect 231394 212548 231400 212560
rect 231268 212520 231400 212548
rect 231268 212508 231274 212520
rect 231394 212508 231400 212520
rect 231452 212508 231458 212560
rect 245028 212492 245056 212644
rect 245010 212440 245016 212492
rect 245068 212440 245074 212492
rect 240686 211080 240692 211132
rect 240744 211120 240750 211132
rect 240870 211120 240876 211132
rect 240744 211092 240876 211120
rect 240744 211080 240750 211092
rect 240870 211080 240876 211092
rect 240928 211080 240934 211132
rect 264330 211080 264336 211132
rect 264388 211120 264394 211132
rect 264514 211120 264520 211132
rect 264388 211092 264520 211120
rect 264388 211080 264394 211092
rect 264514 211080 264520 211092
rect 264572 211080 264578 211132
rect 293126 211080 293132 211132
rect 293184 211120 293190 211132
rect 293310 211120 293316 211132
rect 293184 211092 293316 211120
rect 293184 211080 293190 211092
rect 293310 211080 293316 211092
rect 293368 211080 293374 211132
rect 294598 211080 294604 211132
rect 294656 211120 294662 211132
rect 294782 211120 294788 211132
rect 294656 211092 294788 211120
rect 294656 211080 294662 211092
rect 294782 211080 294788 211092
rect 294840 211080 294846 211132
rect 295886 211080 295892 211132
rect 295944 211120 295950 211132
rect 296070 211120 296076 211132
rect 295944 211092 296076 211120
rect 295944 211080 295950 211092
rect 296070 211080 296076 211092
rect 296128 211080 296134 211132
rect 340046 211120 340052 211132
rect 340007 211092 340052 211120
rect 340046 211080 340052 211092
rect 340104 211080 340110 211132
rect 246390 209828 246396 209840
rect 246351 209800 246396 209828
rect 246390 209788 246396 209800
rect 246448 209788 246454 209840
rect 319622 209828 319628 209840
rect 319583 209800 319628 209828
rect 319622 209788 319628 209800
rect 319680 209788 319686 209840
rect 321094 209828 321100 209840
rect 321055 209800 321100 209828
rect 321094 209788 321100 209800
rect 321152 209788 321158 209840
rect 322106 209828 322112 209840
rect 322067 209800 322112 209828
rect 322106 209788 322112 209800
rect 322164 209788 322170 209840
rect 335814 209760 335820 209772
rect 335775 209732 335820 209760
rect 335814 209720 335820 209732
rect 335872 209720 335878 209772
rect 299014 208496 299020 208548
rect 299072 208496 299078 208548
rect 299032 208412 299060 208496
rect 331766 208428 331772 208480
rect 331824 208428 331830 208480
rect 299014 208360 299020 208412
rect 299072 208360 299078 208412
rect 331784 208400 331812 208428
rect 331858 208400 331864 208412
rect 331784 208372 331864 208400
rect 331858 208360 331864 208372
rect 331916 208360 331922 208412
rect 300302 208332 300308 208344
rect 300263 208304 300308 208332
rect 300302 208292 300308 208304
rect 300360 208292 300366 208344
rect 267182 207748 267188 207800
rect 267240 207748 267246 207800
rect 268654 207748 268660 207800
rect 268712 207748 268718 207800
rect 267200 207664 267228 207748
rect 268672 207664 268700 207748
rect 267182 207612 267188 207664
rect 267240 207612 267246 207664
rect 268654 207612 268660 207664
rect 268712 207612 268718 207664
rect 301590 207000 301596 207052
rect 301648 207040 301654 207052
rect 301777 207043 301835 207049
rect 301777 207040 301789 207043
rect 301648 207012 301789 207040
rect 301648 207000 301654 207012
rect 301777 207009 301789 207012
rect 301823 207009 301835 207043
rect 301777 207003 301835 207009
rect 334618 207000 334624 207052
rect 334676 207040 334682 207052
rect 334676 207012 334721 207040
rect 334676 207000 334682 207012
rect 246390 205640 246396 205692
rect 246448 205640 246454 205692
rect 329009 205683 329067 205689
rect 329009 205649 329021 205683
rect 329055 205680 329067 205683
rect 329098 205680 329104 205692
rect 329055 205652 329104 205680
rect 329055 205649 329067 205652
rect 329009 205643 329067 205649
rect 329098 205640 329104 205652
rect 329156 205640 329162 205692
rect 344094 205640 344100 205692
rect 344152 205680 344158 205692
rect 344278 205680 344284 205692
rect 344152 205652 344284 205680
rect 344152 205640 344158 205652
rect 344278 205640 344284 205652
rect 344336 205640 344342 205692
rect 246408 205544 246436 205640
rect 262858 205572 262864 205624
rect 262916 205612 262922 205624
rect 263042 205612 263048 205624
rect 262916 205584 263048 205612
rect 262916 205572 262922 205584
rect 263042 205572 263048 205584
rect 263100 205572 263106 205624
rect 330573 205615 330631 205621
rect 330573 205581 330585 205615
rect 330619 205612 330631 205615
rect 330754 205612 330760 205624
rect 330619 205584 330760 205612
rect 330619 205581 330631 205584
rect 330573 205575 330631 205581
rect 330754 205572 330760 205584
rect 330812 205572 330818 205624
rect 246482 205544 246488 205556
rect 246408 205516 246488 205544
rect 246482 205504 246488 205516
rect 246540 205504 246546 205556
rect 340049 204935 340107 204941
rect 340049 204901 340061 204935
rect 340095 204932 340107 204935
rect 340230 204932 340236 204944
rect 340095 204904 340236 204932
rect 340095 204901 340107 204904
rect 340049 204895 340107 204901
rect 340230 204892 340236 204904
rect 340288 204892 340294 204944
rect 261570 203600 261576 203652
rect 261628 203640 261634 203652
rect 261662 203640 261668 203652
rect 261628 203612 261668 203640
rect 261628 203600 261634 203612
rect 261662 203600 261668 203612
rect 261720 203600 261726 203652
rect 335817 203575 335875 203581
rect 335817 203541 335829 203575
rect 335863 203572 335875 203575
rect 336090 203572 336096 203584
rect 335863 203544 336096 203572
rect 335863 203541 335875 203544
rect 335817 203535 335875 203541
rect 336090 203532 336096 203544
rect 336148 203532 336154 203584
rect 244550 202920 244556 202972
rect 244608 202920 244614 202972
rect 257154 202960 257160 202972
rect 257080 202932 257160 202960
rect 100662 202852 100668 202904
rect 100720 202892 100726 202904
rect 100846 202892 100852 202904
rect 100720 202864 100852 202892
rect 100720 202852 100726 202864
rect 100846 202852 100852 202864
rect 100904 202852 100910 202904
rect 232314 202852 232320 202904
rect 232372 202892 232378 202904
rect 232590 202892 232596 202904
rect 232372 202864 232596 202892
rect 232372 202852 232378 202864
rect 232590 202852 232596 202864
rect 232648 202852 232654 202904
rect 238018 202852 238024 202904
rect 238076 202892 238082 202904
rect 238110 202892 238116 202904
rect 238076 202864 238116 202892
rect 238076 202852 238082 202864
rect 238110 202852 238116 202864
rect 238168 202852 238174 202904
rect 244458 202892 244464 202904
rect 244419 202864 244464 202892
rect 244458 202852 244464 202864
rect 244516 202852 244522 202904
rect 244568 202836 244596 202920
rect 257080 202904 257108 202932
rect 257154 202920 257160 202932
rect 257212 202920 257218 202972
rect 253014 202852 253020 202904
rect 253072 202892 253078 202904
rect 253106 202892 253112 202904
rect 253072 202864 253112 202892
rect 253072 202852 253078 202864
rect 253106 202852 253112 202864
rect 253164 202852 253170 202904
rect 257062 202852 257068 202904
rect 257120 202852 257126 202904
rect 258718 202852 258724 202904
rect 258776 202892 258782 202904
rect 258810 202892 258816 202904
rect 258776 202864 258816 202892
rect 258776 202852 258782 202864
rect 258810 202852 258816 202864
rect 258868 202852 258874 202904
rect 260282 202852 260288 202904
rect 260340 202892 260346 202904
rect 260374 202892 260380 202904
rect 260340 202864 260380 202892
rect 260340 202852 260346 202864
rect 260374 202852 260380 202864
rect 260432 202852 260438 202904
rect 244550 202784 244556 202836
rect 244608 202784 244614 202836
rect 244458 201532 244464 201544
rect 244419 201504 244464 201532
rect 244458 201492 244464 201504
rect 244516 201492 244522 201544
rect 107470 201424 107476 201476
rect 107528 201464 107534 201476
rect 107654 201464 107660 201476
rect 107528 201436 107660 201464
rect 107528 201424 107534 201436
rect 107654 201424 107660 201436
rect 107712 201424 107718 201476
rect 264330 201424 264336 201476
rect 264388 201464 264394 201476
rect 264514 201464 264520 201476
rect 264388 201436 264520 201464
rect 264388 201424 264394 201436
rect 264514 201424 264520 201436
rect 264572 201424 264578 201476
rect 293126 201424 293132 201476
rect 293184 201464 293190 201476
rect 293310 201464 293316 201476
rect 293184 201436 293316 201464
rect 293184 201424 293190 201436
rect 293310 201424 293316 201436
rect 293368 201424 293374 201476
rect 345382 201424 345388 201476
rect 345440 201464 345446 201476
rect 345566 201464 345572 201476
rect 345440 201436 345572 201464
rect 345440 201424 345446 201436
rect 345566 201424 345572 201436
rect 345624 201424 345630 201476
rect 326246 200172 326252 200184
rect 326207 200144 326252 200172
rect 326246 200132 326252 200144
rect 326304 200132 326310 200184
rect 319622 200104 319628 200116
rect 319583 200076 319628 200104
rect 319622 200064 319628 200076
rect 319680 200064 319686 200116
rect 321094 200104 321100 200116
rect 321055 200076 321100 200104
rect 321094 200064 321100 200076
rect 321152 200064 321158 200116
rect 322201 200107 322259 200113
rect 322201 200073 322213 200107
rect 322247 200104 322259 200107
rect 322290 200104 322296 200116
rect 322247 200076 322296 200104
rect 322247 200073 322259 200076
rect 322201 200067 322259 200073
rect 322290 200064 322296 200076
rect 322348 200064 322354 200116
rect 300302 198744 300308 198756
rect 300263 198716 300308 198744
rect 300302 198704 300308 198716
rect 300360 198704 300366 198756
rect 299014 198676 299020 198688
rect 298975 198648 299020 198676
rect 299014 198636 299020 198648
rect 299072 198636 299078 198688
rect 301774 197276 301780 197328
rect 301832 197276 301838 197328
rect 329009 197319 329067 197325
rect 329009 197285 329021 197319
rect 329055 197316 329067 197319
rect 329098 197316 329104 197328
rect 329055 197288 329104 197316
rect 329055 197285 329067 197288
rect 329009 197279 329067 197285
rect 329098 197276 329104 197288
rect 329156 197276 329162 197328
rect 331858 197276 331864 197328
rect 331916 197316 331922 197328
rect 332042 197316 332048 197328
rect 331916 197288 332048 197316
rect 331916 197276 331922 197288
rect 332042 197276 332048 197288
rect 332100 197276 332106 197328
rect 334618 197316 334624 197328
rect 334579 197288 334624 197316
rect 334618 197276 334624 197288
rect 334676 197276 334682 197328
rect 301792 197189 301820 197276
rect 301777 197183 301835 197189
rect 301777 197149 301789 197183
rect 301823 197149 301835 197183
rect 301777 197143 301835 197149
rect 326246 196052 326252 196104
rect 326304 196052 326310 196104
rect 232774 196024 232780 196036
rect 232700 195996 232780 196024
rect 232700 195968 232728 195996
rect 232774 195984 232780 195996
rect 232832 195984 232838 196036
rect 326264 195968 326292 196052
rect 232682 195916 232688 195968
rect 232740 195916 232746 195968
rect 326246 195916 326252 195968
rect 326304 195916 326310 195968
rect 341518 195916 341524 195968
rect 341576 195956 341582 195968
rect 341702 195956 341708 195968
rect 341576 195928 341708 195956
rect 341576 195916 341582 195928
rect 341702 195916 341708 195928
rect 341760 195916 341766 195968
rect 244921 195279 244979 195285
rect 244921 195245 244933 195279
rect 244967 195276 244979 195279
rect 245010 195276 245016 195288
rect 244967 195248 245016 195276
rect 244967 195245 244979 195248
rect 244921 195239 244979 195245
rect 245010 195236 245016 195248
rect 245068 195236 245074 195288
rect 2774 194284 2780 194336
rect 2832 194324 2838 194336
rect 5074 194324 5080 194336
rect 2832 194296 5080 194324
rect 2832 194284 2838 194296
rect 5074 194284 5080 194296
rect 5132 194284 5138 194336
rect 231210 193196 231216 193248
rect 231268 193236 231274 193248
rect 231394 193236 231400 193248
rect 231268 193208 231400 193236
rect 231268 193196 231274 193208
rect 231394 193196 231400 193208
rect 231452 193196 231458 193248
rect 232314 193196 232320 193248
rect 232372 193236 232378 193248
rect 232406 193236 232412 193248
rect 232372 193208 232412 193236
rect 232372 193196 232378 193208
rect 232406 193196 232412 193208
rect 232464 193196 232470 193248
rect 246390 193196 246396 193248
rect 246448 193236 246454 193248
rect 246574 193236 246580 193248
rect 246448 193208 246580 193236
rect 246448 193196 246454 193208
rect 246574 193196 246580 193208
rect 246632 193196 246638 193248
rect 333054 193196 333060 193248
rect 333112 193236 333118 193248
rect 333146 193236 333152 193248
rect 333112 193208 333152 193236
rect 333112 193196 333118 193208
rect 333146 193196 333152 193208
rect 333204 193196 333210 193248
rect 253014 191836 253020 191888
rect 253072 191876 253078 191888
rect 253106 191876 253112 191888
rect 253072 191848 253112 191876
rect 253072 191836 253078 191848
rect 253106 191836 253112 191848
rect 253164 191836 253170 191888
rect 258810 191836 258816 191888
rect 258868 191876 258874 191888
rect 258902 191876 258908 191888
rect 258868 191848 258908 191876
rect 258868 191836 258874 191848
rect 258902 191836 258908 191848
rect 258960 191836 258966 191888
rect 232130 191768 232136 191820
rect 232188 191808 232194 191820
rect 232406 191808 232412 191820
rect 232188 191780 232412 191808
rect 232188 191768 232194 191780
rect 232406 191768 232412 191780
rect 232464 191768 232470 191820
rect 240686 191768 240692 191820
rect 240744 191768 240750 191820
rect 260190 191808 260196 191820
rect 260151 191780 260196 191808
rect 260190 191768 260196 191780
rect 260248 191768 260254 191820
rect 264330 191768 264336 191820
rect 264388 191808 264394 191820
rect 264514 191808 264520 191820
rect 264388 191780 264520 191808
rect 264388 191768 264394 191780
rect 264514 191768 264520 191780
rect 264572 191768 264578 191820
rect 265618 191768 265624 191820
rect 265676 191808 265682 191820
rect 265802 191808 265808 191820
rect 265676 191780 265808 191808
rect 265676 191768 265682 191780
rect 265802 191768 265808 191780
rect 265860 191768 265866 191820
rect 293126 191768 293132 191820
rect 293184 191808 293190 191820
rect 293310 191808 293316 191820
rect 293184 191780 293316 191808
rect 293184 191768 293190 191780
rect 293310 191768 293316 191780
rect 293368 191768 293374 191820
rect 294598 191768 294604 191820
rect 294656 191808 294662 191820
rect 294782 191808 294788 191820
rect 294656 191780 294788 191808
rect 294656 191768 294662 191780
rect 294782 191768 294788 191780
rect 294840 191768 294846 191820
rect 295886 191768 295892 191820
rect 295944 191808 295950 191820
rect 296070 191808 296076 191820
rect 295944 191780 296076 191808
rect 295944 191768 295950 191780
rect 296070 191768 296076 191780
rect 296128 191768 296134 191820
rect 333054 191768 333060 191820
rect 333112 191808 333118 191820
rect 333146 191808 333152 191820
rect 333112 191780 333152 191808
rect 333112 191768 333118 191780
rect 333146 191768 333152 191780
rect 333204 191768 333210 191820
rect 240704 191740 240732 191768
rect 240870 191740 240876 191752
rect 240704 191712 240876 191740
rect 240870 191700 240876 191712
rect 240928 191700 240934 191752
rect 319622 190516 319628 190528
rect 319583 190488 319628 190516
rect 319622 190476 319628 190488
rect 319680 190476 319686 190528
rect 321094 190516 321100 190528
rect 321055 190488 321100 190516
rect 321094 190476 321100 190488
rect 321152 190476 321158 190528
rect 322198 190516 322204 190528
rect 322159 190488 322204 190516
rect 322198 190476 322204 190488
rect 322256 190476 322262 190528
rect 261478 190448 261484 190460
rect 261439 190420 261484 190448
rect 261478 190408 261484 190420
rect 261536 190408 261542 190460
rect 263042 190448 263048 190460
rect 263003 190420 263048 190448
rect 263042 190408 263048 190420
rect 263100 190408 263106 190460
rect 333238 190408 333244 190460
rect 333296 190448 333302 190460
rect 333330 190448 333336 190460
rect 333296 190420 333336 190448
rect 333296 190408 333302 190420
rect 333330 190408 333336 190420
rect 333388 190408 333394 190460
rect 335814 190448 335820 190460
rect 335775 190420 335820 190448
rect 335814 190408 335820 190420
rect 335872 190408 335878 190460
rect 244182 189456 244188 189508
rect 244240 189496 244246 189508
rect 244369 189499 244427 189505
rect 244369 189496 244381 189499
rect 244240 189468 244381 189496
rect 244240 189456 244246 189468
rect 244369 189465 244381 189468
rect 244415 189465 244427 189499
rect 244369 189459 244427 189465
rect 299014 189088 299020 189100
rect 298975 189060 299020 189088
rect 299014 189048 299020 189060
rect 299072 189048 299078 189100
rect 300302 189020 300308 189032
rect 300263 188992 300308 189020
rect 300302 188980 300308 188992
rect 300360 188980 300366 189032
rect 301774 187728 301780 187740
rect 301735 187700 301780 187728
rect 301774 187688 301780 187700
rect 301832 187688 301838 187740
rect 329006 187728 329012 187740
rect 328967 187700 329012 187728
rect 329006 187688 329012 187700
rect 329064 187688 329070 187740
rect 330570 187728 330576 187740
rect 330531 187700 330576 187728
rect 330570 187688 330576 187700
rect 330628 187688 330634 187740
rect 334618 187728 334624 187740
rect 334579 187700 334624 187728
rect 334618 187688 334624 187700
rect 334676 187688 334682 187740
rect 257154 186436 257160 186448
rect 257080 186408 257160 186436
rect 257080 186312 257108 186408
rect 257154 186396 257160 186408
rect 257212 186396 257218 186448
rect 258902 186328 258908 186380
rect 258960 186328 258966 186380
rect 257062 186260 257068 186312
rect 257120 186260 257126 186312
rect 258920 186244 258948 186328
rect 258902 186192 258908 186244
rect 258960 186192 258966 186244
rect 333146 183920 333152 183932
rect 333107 183892 333152 183920
rect 333146 183880 333152 183892
rect 333204 183880 333210 183932
rect 345382 183648 345388 183660
rect 345308 183620 345388 183648
rect 345308 183592 345336 183620
rect 345382 183608 345388 183620
rect 345440 183608 345446 183660
rect 100662 183540 100668 183592
rect 100720 183580 100726 183592
rect 100846 183580 100852 183592
rect 100720 183552 100852 183580
rect 100720 183540 100726 183552
rect 100846 183540 100852 183552
rect 100904 183540 100910 183592
rect 238018 183540 238024 183592
rect 238076 183580 238082 183592
rect 238110 183580 238116 183592
rect 238076 183552 238116 183580
rect 238076 183540 238082 183552
rect 238110 183540 238116 183552
rect 238168 183540 238174 183592
rect 244921 183583 244979 183589
rect 244921 183549 244933 183583
rect 244967 183580 244979 183583
rect 245010 183580 245016 183592
rect 244967 183552 245016 183580
rect 244967 183549 244979 183552
rect 244921 183543 244979 183549
rect 245010 183540 245016 183552
rect 245068 183540 245074 183592
rect 341610 183540 341616 183592
rect 341668 183580 341674 183592
rect 341702 183580 341708 183592
rect 341668 183552 341708 183580
rect 341668 183540 341674 183552
rect 341702 183540 341708 183552
rect 341760 183540 341766 183592
rect 345290 183540 345296 183592
rect 345348 183540 345354 183592
rect 260193 183515 260251 183521
rect 260193 183481 260205 183515
rect 260239 183512 260251 183515
rect 260282 183512 260288 183524
rect 260239 183484 260288 183512
rect 260239 183481 260251 183484
rect 260193 183475 260251 183481
rect 260282 183472 260288 183484
rect 260340 183472 260346 183524
rect 107470 182112 107476 182164
rect 107528 182152 107534 182164
rect 107654 182152 107660 182164
rect 107528 182124 107660 182152
rect 107528 182112 107534 182124
rect 107654 182112 107660 182124
rect 107712 182112 107718 182164
rect 232038 182112 232044 182164
rect 232096 182112 232102 182164
rect 232314 182152 232320 182164
rect 232275 182124 232320 182152
rect 232314 182112 232320 182124
rect 232372 182112 232378 182164
rect 260282 182152 260288 182164
rect 260243 182124 260288 182152
rect 260282 182112 260288 182124
rect 260340 182112 260346 182164
rect 261478 182152 261484 182164
rect 261439 182124 261484 182152
rect 261478 182112 261484 182124
rect 261536 182112 261542 182164
rect 293126 182112 293132 182164
rect 293184 182152 293190 182164
rect 293310 182152 293316 182164
rect 293184 182124 293316 182152
rect 293184 182112 293190 182124
rect 293310 182112 293316 182124
rect 293368 182112 293374 182164
rect 231946 182044 231952 182096
rect 232004 182084 232010 182096
rect 232056 182084 232084 182112
rect 333146 182084 333152 182096
rect 232004 182056 232084 182084
rect 333107 182056 333152 182084
rect 232004 182044 232010 182056
rect 333146 182044 333152 182056
rect 333204 182044 333210 182096
rect 263042 180820 263048 180872
rect 263100 180860 263106 180872
rect 334529 180863 334587 180869
rect 263100 180832 263145 180860
rect 263100 180820 263106 180832
rect 334529 180829 334541 180863
rect 334575 180860 334587 180863
rect 334618 180860 334624 180872
rect 334575 180832 334624 180860
rect 334575 180829 334587 180832
rect 334529 180823 334587 180829
rect 334618 180820 334624 180832
rect 334676 180820 334682 180872
rect 335814 180860 335820 180872
rect 335775 180832 335820 180860
rect 335814 180820 335820 180832
rect 335872 180820 335878 180872
rect 264514 180792 264520 180804
rect 264475 180764 264520 180792
rect 264514 180752 264520 180764
rect 264572 180752 264578 180804
rect 265802 180792 265808 180804
rect 265763 180764 265808 180792
rect 265802 180752 265808 180764
rect 265860 180752 265866 180804
rect 293126 180792 293132 180804
rect 293087 180764 293132 180792
rect 293126 180752 293132 180764
rect 293184 180752 293190 180804
rect 319622 180792 319628 180804
rect 319583 180764 319628 180792
rect 319622 180752 319628 180764
rect 319680 180752 319686 180804
rect 321094 180792 321100 180804
rect 321055 180764 321100 180792
rect 321094 180752 321100 180764
rect 321152 180752 321158 180804
rect 2774 179664 2780 179716
rect 2832 179704 2838 179716
rect 4982 179704 4988 179716
rect 2832 179676 4988 179704
rect 2832 179664 2838 179676
rect 4982 179664 4988 179676
rect 5040 179664 5046 179716
rect 301774 179596 301780 179648
rect 301832 179596 301838 179648
rect 301792 179512 301820 179596
rect 301774 179460 301780 179512
rect 301832 179460 301838 179512
rect 334526 179500 334532 179512
rect 334487 179472 334532 179500
rect 334526 179460 334532 179472
rect 334584 179460 334590 179512
rect 298922 179392 298928 179444
rect 298980 179432 298986 179444
rect 299014 179432 299020 179444
rect 298980 179404 299020 179432
rect 298980 179392 298986 179404
rect 299014 179392 299020 179404
rect 299072 179392 299078 179444
rect 300302 179432 300308 179444
rect 300263 179404 300308 179432
rect 300302 179392 300308 179404
rect 300360 179392 300366 179444
rect 329006 179324 329012 179376
rect 329064 179364 329070 179376
rect 329098 179364 329104 179376
rect 329064 179336 329104 179364
rect 329064 179324 329070 179336
rect 329098 179324 329104 179336
rect 329156 179324 329162 179376
rect 334526 179364 334532 179376
rect 334487 179336 334532 179364
rect 334526 179324 334532 179336
rect 334584 179324 334590 179376
rect 340046 178780 340052 178832
rect 340104 178780 340110 178832
rect 340064 178752 340092 178780
rect 340138 178752 340144 178764
rect 340064 178724 340144 178752
rect 340138 178712 340144 178724
rect 340196 178712 340202 178764
rect 331858 178032 331864 178084
rect 331916 178072 331922 178084
rect 332042 178072 332048 178084
rect 331916 178044 332048 178072
rect 331916 178032 331922 178044
rect 332042 178032 332048 178044
rect 332100 178032 332106 178084
rect 301774 178004 301780 178016
rect 301735 177976 301780 178004
rect 301774 177964 301780 177976
rect 301832 177964 301838 178016
rect 232682 176604 232688 176656
rect 232740 176604 232746 176656
rect 232700 176520 232728 176604
rect 232682 176468 232688 176520
rect 232740 176468 232746 176520
rect 231210 173884 231216 173936
rect 231268 173924 231274 173936
rect 231394 173924 231400 173936
rect 231268 173896 231400 173924
rect 231268 173884 231274 173896
rect 231394 173884 231400 173896
rect 231452 173884 231458 173936
rect 244369 173927 244427 173933
rect 244369 173893 244381 173927
rect 244415 173924 244427 173927
rect 244458 173924 244464 173936
rect 244415 173896 244464 173924
rect 244415 173893 244427 173896
rect 244369 173887 244427 173893
rect 244458 173884 244464 173896
rect 244516 173884 244522 173936
rect 244918 173884 244924 173936
rect 244976 173924 244982 173936
rect 245102 173924 245108 173936
rect 244976 173896 245108 173924
rect 244976 173884 244982 173896
rect 245102 173884 245108 173896
rect 245160 173884 245166 173936
rect 245838 173884 245844 173936
rect 245896 173924 245902 173936
rect 246022 173924 246028 173936
rect 245896 173896 246028 173924
rect 245896 173884 245902 173896
rect 246022 173884 246028 173896
rect 246080 173884 246086 173936
rect 246390 173884 246396 173936
rect 246448 173924 246454 173936
rect 246574 173924 246580 173936
rect 246448 173896 246580 173924
rect 246448 173884 246454 173896
rect 246574 173884 246580 173896
rect 246632 173884 246638 173936
rect 333238 173884 333244 173936
rect 333296 173884 333302 173936
rect 335814 173884 335820 173936
rect 335872 173884 335878 173936
rect 345290 173884 345296 173936
rect 345348 173924 345354 173936
rect 345382 173924 345388 173936
rect 345348 173896 345388 173924
rect 345348 173884 345354 173896
rect 345382 173884 345388 173896
rect 345440 173884 345446 173936
rect 260282 173856 260288 173868
rect 260243 173828 260288 173856
rect 260282 173816 260288 173828
rect 260340 173816 260346 173868
rect 333256 173788 333284 173884
rect 333330 173788 333336 173800
rect 333256 173760 333336 173788
rect 333330 173748 333336 173760
rect 333388 173748 333394 173800
rect 335832 173788 335860 173884
rect 335906 173788 335912 173800
rect 335832 173760 335912 173788
rect 335906 173748 335912 173760
rect 335964 173748 335970 173800
rect 232317 172567 232375 172573
rect 232317 172533 232329 172567
rect 232363 172564 232375 172567
rect 232406 172564 232412 172576
rect 232363 172536 232412 172564
rect 232363 172533 232375 172536
rect 232317 172527 232375 172533
rect 232406 172524 232412 172536
rect 232464 172524 232470 172576
rect 252922 172524 252928 172576
rect 252980 172564 252986 172576
rect 253014 172564 253020 172576
rect 252980 172536 253020 172564
rect 252980 172524 252986 172536
rect 253014 172524 253020 172536
rect 253072 172524 253078 172576
rect 256970 172524 256976 172576
rect 257028 172564 257034 172576
rect 257062 172564 257068 172576
rect 257028 172536 257068 172564
rect 257028 172524 257034 172536
rect 257062 172524 257068 172536
rect 257120 172524 257126 172576
rect 258810 172524 258816 172576
rect 258868 172564 258874 172576
rect 258902 172564 258908 172576
rect 258868 172536 258908 172564
rect 258868 172524 258874 172536
rect 258902 172524 258908 172536
rect 258960 172524 258966 172576
rect 240686 172456 240692 172508
rect 240744 172496 240750 172508
rect 240870 172496 240876 172508
rect 240744 172468 240876 172496
rect 240744 172456 240750 172468
rect 240870 172456 240876 172468
rect 240928 172456 240934 172508
rect 294782 171232 294788 171284
rect 294840 171232 294846 171284
rect 296070 171232 296076 171284
rect 296128 171232 296134 171284
rect 294800 171148 294828 171232
rect 296088 171148 296116 171232
rect 322290 171164 322296 171216
rect 322348 171164 322354 171216
rect 264514 171136 264520 171148
rect 264475 171108 264520 171136
rect 264514 171096 264520 171108
rect 264572 171096 264578 171148
rect 265802 171136 265808 171148
rect 265763 171108 265808 171136
rect 265802 171096 265808 171108
rect 265860 171096 265866 171148
rect 293129 171139 293187 171145
rect 293129 171105 293141 171139
rect 293175 171136 293187 171139
rect 293310 171136 293316 171148
rect 293175 171108 293316 171136
rect 293175 171105 293187 171108
rect 293129 171099 293187 171105
rect 293310 171096 293316 171108
rect 293368 171096 293374 171148
rect 294782 171096 294788 171148
rect 294840 171096 294846 171148
rect 296070 171096 296076 171148
rect 296128 171096 296134 171148
rect 319622 171136 319628 171148
rect 319583 171108 319628 171136
rect 319622 171096 319628 171108
rect 319680 171096 319686 171148
rect 321094 171136 321100 171148
rect 321055 171108 321100 171136
rect 321094 171096 321100 171108
rect 321152 171096 321158 171148
rect 322308 171136 322336 171164
rect 322382 171136 322388 171148
rect 322308 171108 322388 171136
rect 322382 171096 322388 171108
rect 322440 171096 322446 171148
rect 334526 171068 334532 171080
rect 334487 171040 334532 171068
rect 334526 171028 334532 171040
rect 334584 171028 334590 171080
rect 331769 169847 331827 169853
rect 331769 169813 331781 169847
rect 331815 169844 331827 169847
rect 331858 169844 331864 169856
rect 331815 169816 331864 169844
rect 331815 169813 331827 169816
rect 331769 169807 331827 169813
rect 331858 169804 331864 169816
rect 331916 169804 331922 169856
rect 299014 169708 299020 169720
rect 298975 169680 299020 169708
rect 299014 169668 299020 169680
rect 299072 169668 299078 169720
rect 300302 169708 300308 169720
rect 300263 169680 300308 169708
rect 300302 169668 300308 169680
rect 300360 169668 300366 169720
rect 326338 169708 326344 169720
rect 326299 169680 326344 169708
rect 326338 169668 326344 169680
rect 326396 169668 326402 169720
rect 340138 169056 340144 169108
rect 340196 169096 340202 169108
rect 340322 169096 340328 169108
rect 340196 169068 340328 169096
rect 340196 169056 340202 169068
rect 340322 169056 340328 169068
rect 340380 169056 340386 169108
rect 301774 168416 301780 168428
rect 301735 168388 301780 168416
rect 301774 168376 301780 168388
rect 301832 168376 301838 168428
rect 331766 168416 331772 168428
rect 331727 168388 331772 168416
rect 331766 168376 331772 168388
rect 331824 168376 331830 168428
rect 231946 167628 231952 167680
rect 232004 167668 232010 167680
rect 232130 167668 232136 167680
rect 232004 167640 232136 167668
rect 232004 167628 232010 167640
rect 232130 167628 232136 167640
rect 232188 167628 232194 167680
rect 322382 167084 322388 167136
rect 322440 167084 322446 167136
rect 232406 167056 232412 167068
rect 232332 167028 232412 167056
rect 232332 167000 232360 167028
rect 232406 167016 232412 167028
rect 232464 167016 232470 167068
rect 232314 166948 232320 167000
rect 232372 166948 232378 167000
rect 322290 166880 322296 166932
rect 322348 166920 322354 166932
rect 322400 166920 322428 167084
rect 322348 166892 322428 166920
rect 322348 166880 322354 166892
rect 335906 166268 335912 166320
rect 335964 166308 335970 166320
rect 336090 166308 336096 166320
rect 335964 166280 336096 166308
rect 335964 166268 335970 166280
rect 336090 166268 336096 166280
rect 336148 166268 336154 166320
rect 261662 164336 261668 164348
rect 261588 164308 261668 164336
rect 261588 164280 261616 164308
rect 261662 164296 261668 164308
rect 261720 164296 261726 164348
rect 252922 164228 252928 164280
rect 252980 164268 252986 164280
rect 253014 164268 253020 164280
rect 252980 164240 253020 164268
rect 252980 164228 252986 164240
rect 253014 164228 253020 164240
rect 253072 164228 253078 164280
rect 256970 164228 256976 164280
rect 257028 164268 257034 164280
rect 257062 164268 257068 164280
rect 257028 164240 257068 164268
rect 257028 164228 257034 164240
rect 257062 164228 257068 164240
rect 257120 164228 257126 164280
rect 261570 164228 261576 164280
rect 261628 164228 261634 164280
rect 244182 164160 244188 164212
rect 244240 164200 244246 164212
rect 244366 164200 244372 164212
rect 244240 164172 244372 164200
rect 244240 164160 244246 164172
rect 244366 164160 244372 164172
rect 244424 164160 244430 164212
rect 340046 164160 340052 164212
rect 340104 164200 340110 164212
rect 340138 164200 340144 164212
rect 340104 164172 340144 164200
rect 340104 164160 340110 164172
rect 340138 164160 340144 164172
rect 340196 164160 340202 164212
rect 345382 164160 345388 164212
rect 345440 164200 345446 164212
rect 345566 164200 345572 164212
rect 345440 164172 345572 164200
rect 345440 164160 345446 164172
rect 345566 164160 345572 164172
rect 345624 164160 345630 164212
rect 107470 162840 107476 162852
rect 107431 162812 107476 162840
rect 107470 162800 107476 162812
rect 107528 162800 107534 162852
rect 232038 162800 232044 162852
rect 232096 162840 232102 162852
rect 232130 162840 232136 162852
rect 232096 162812 232136 162840
rect 232096 162800 232102 162812
rect 232130 162800 232136 162812
rect 232188 162800 232194 162852
rect 232314 162800 232320 162852
rect 232372 162840 232378 162852
rect 232590 162840 232596 162852
rect 232372 162812 232596 162840
rect 232372 162800 232378 162812
rect 232590 162800 232596 162812
rect 232648 162800 232654 162852
rect 261570 162800 261576 162852
rect 261628 162840 261634 162852
rect 261662 162840 261668 162852
rect 261628 162812 261668 162840
rect 261628 162800 261634 162812
rect 261662 162800 261668 162812
rect 261720 162800 261726 162852
rect 329006 161440 329012 161492
rect 329064 161480 329070 161492
rect 329098 161480 329104 161492
rect 329064 161452 329104 161480
rect 329064 161440 329070 161452
rect 329098 161440 329104 161452
rect 329156 161440 329162 161492
rect 232590 161412 232596 161424
rect 232551 161384 232596 161412
rect 232590 161372 232596 161384
rect 232648 161372 232654 161424
rect 253014 161412 253020 161424
rect 252975 161384 253020 161412
rect 253014 161372 253020 161384
rect 253072 161372 253078 161424
rect 257062 161412 257068 161424
rect 257023 161384 257068 161412
rect 257062 161372 257068 161384
rect 257120 161372 257126 161424
rect 293310 161412 293316 161424
rect 293271 161384 293316 161412
rect 293310 161372 293316 161384
rect 293368 161372 293374 161424
rect 319622 161412 319628 161424
rect 319583 161384 319628 161412
rect 319622 161372 319628 161384
rect 319680 161372 319686 161424
rect 321094 161412 321100 161424
rect 321055 161384 321100 161412
rect 321094 161372 321100 161384
rect 321152 161372 321158 161424
rect 326341 161347 326399 161353
rect 326341 161313 326353 161347
rect 326387 161344 326399 161347
rect 326430 161344 326436 161356
rect 326387 161316 326436 161344
rect 326387 161313 326399 161316
rect 326341 161307 326399 161313
rect 326430 161304 326436 161316
rect 326488 161304 326494 161356
rect 301866 160352 301872 160404
rect 301924 160352 301930 160404
rect 301884 160132 301912 160352
rect 299014 160120 299020 160132
rect 298975 160092 299020 160120
rect 299014 160080 299020 160092
rect 299072 160080 299078 160132
rect 300302 160120 300308 160132
rect 300263 160092 300308 160120
rect 300302 160080 300308 160092
rect 300360 160080 300366 160132
rect 301774 160080 301780 160132
rect 301832 160080 301838 160132
rect 301866 160080 301872 160132
rect 301924 160080 301930 160132
rect 330478 160080 330484 160132
rect 330536 160120 330542 160132
rect 330570 160120 330576 160132
rect 330536 160092 330576 160120
rect 330536 160080 330542 160092
rect 330570 160080 330576 160092
rect 330628 160080 330634 160132
rect 260374 160012 260380 160064
rect 260432 160012 260438 160064
rect 260282 159944 260288 159996
rect 260340 159984 260346 159996
rect 260392 159984 260420 160012
rect 301792 159996 301820 160080
rect 260340 159956 260420 159984
rect 260340 159944 260346 159956
rect 301774 159944 301780 159996
rect 301832 159944 301838 159996
rect 260282 158692 260288 158704
rect 260243 158664 260288 158692
rect 260282 158652 260288 158664
rect 260340 158652 260346 158704
rect 258810 157428 258816 157480
rect 258868 157428 258874 157480
rect 258828 157344 258856 157428
rect 231210 157292 231216 157344
rect 231268 157292 231274 157344
rect 258810 157292 258816 157344
rect 258868 157292 258874 157344
rect 231228 157208 231256 157292
rect 231210 157156 231216 157208
rect 231268 157156 231274 157208
rect 100662 154504 100668 154556
rect 100720 154544 100726 154556
rect 100846 154544 100852 154556
rect 100720 154516 100852 154544
rect 100720 154504 100726 154516
rect 100846 154504 100852 154516
rect 100904 154504 100910 154556
rect 231210 154504 231216 154556
rect 231268 154544 231274 154556
rect 231394 154544 231400 154556
rect 231268 154516 231400 154544
rect 231268 154504 231274 154516
rect 231394 154504 231400 154516
rect 231452 154504 231458 154556
rect 107470 153252 107476 153264
rect 107431 153224 107476 153252
rect 107470 153212 107476 153224
rect 107528 153212 107534 153264
rect 257246 153212 257252 153264
rect 257304 153212 257310 153264
rect 232041 153187 232099 153193
rect 232041 153153 232053 153187
rect 232087 153184 232099 153187
rect 232130 153184 232136 153196
rect 232087 153156 232136 153184
rect 232087 153153 232099 153156
rect 232041 153147 232099 153153
rect 232130 153144 232136 153156
rect 232188 153144 232194 153196
rect 232590 153184 232596 153196
rect 232551 153156 232596 153184
rect 232590 153144 232596 153156
rect 232648 153144 232654 153196
rect 240686 153144 240692 153196
rect 240744 153184 240750 153196
rect 240870 153184 240876 153196
rect 240744 153156 240876 153184
rect 240744 153144 240750 153156
rect 240870 153144 240876 153156
rect 240928 153144 240934 153196
rect 257264 153128 257292 153212
rect 257246 153076 257252 153128
rect 257304 153076 257310 153128
rect 294782 151920 294788 151972
rect 294840 151920 294846 151972
rect 296070 151920 296076 151972
rect 296128 151920 296134 151972
rect 294800 151836 294828 151920
rect 296088 151836 296116 151920
rect 253014 151824 253020 151836
rect 252975 151796 253020 151824
rect 253014 151784 253020 151796
rect 253072 151784 253078 151836
rect 257065 151827 257123 151833
rect 257065 151793 257077 151827
rect 257111 151824 257123 151827
rect 257338 151824 257344 151836
rect 257111 151796 257344 151824
rect 257111 151793 257123 151796
rect 257065 151787 257123 151793
rect 257338 151784 257344 151796
rect 257396 151784 257402 151836
rect 293310 151824 293316 151836
rect 293271 151796 293316 151824
rect 293310 151784 293316 151796
rect 293368 151784 293374 151836
rect 294782 151784 294788 151836
rect 294840 151784 294846 151836
rect 296070 151784 296076 151836
rect 296128 151784 296134 151836
rect 319622 151824 319628 151836
rect 319583 151796 319628 151824
rect 319622 151784 319628 151796
rect 319680 151784 319686 151836
rect 321094 151824 321100 151836
rect 321055 151796 321100 151824
rect 321094 151784 321100 151796
rect 321152 151784 321158 151836
rect 333238 151784 333244 151836
rect 333296 151824 333302 151836
rect 333330 151824 333336 151836
rect 333296 151796 333336 151824
rect 333296 151784 333302 151796
rect 333330 151784 333336 151796
rect 333388 151784 333394 151836
rect 264514 151756 264520 151768
rect 264475 151728 264520 151756
rect 264514 151716 264520 151728
rect 264572 151716 264578 151768
rect 322290 151716 322296 151768
rect 322348 151756 322354 151768
rect 322382 151756 322388 151768
rect 322348 151728 322388 151756
rect 322348 151716 322354 151728
rect 322382 151716 322388 151728
rect 322440 151716 322446 151768
rect 331766 151756 331772 151768
rect 331727 151728 331772 151756
rect 331766 151716 331772 151728
rect 331824 151716 331830 151768
rect 334526 151756 334532 151768
rect 334487 151728 334532 151756
rect 334526 151716 334532 151728
rect 334584 151716 334590 151768
rect 253014 151688 253020 151700
rect 252975 151660 253020 151688
rect 253014 151648 253020 151660
rect 253072 151648 253078 151700
rect 2774 151308 2780 151360
rect 2832 151348 2838 151360
rect 4890 151348 4896 151360
rect 2832 151320 4896 151348
rect 2832 151308 2838 151320
rect 4890 151308 4896 151320
rect 4948 151308 4954 151360
rect 296070 150396 296076 150408
rect 296031 150368 296076 150396
rect 296070 150356 296076 150368
rect 296128 150356 296134 150408
rect 330478 150396 330484 150408
rect 330439 150368 330484 150396
rect 330478 150356 330484 150368
rect 330536 150356 330542 150408
rect 301501 150263 301559 150269
rect 301501 150229 301513 150263
rect 301547 150260 301559 150263
rect 301774 150260 301780 150272
rect 301547 150232 301780 150260
rect 301547 150229 301559 150232
rect 301501 150223 301559 150229
rect 301774 150220 301780 150232
rect 301832 150220 301838 150272
rect 260282 149104 260288 149116
rect 260243 149076 260288 149104
rect 260282 149064 260288 149076
rect 260340 149064 260346 149116
rect 244458 147744 244464 147756
rect 244384 147716 244464 147744
rect 244384 147620 244412 147716
rect 244458 147704 244464 147716
rect 244516 147704 244522 147756
rect 244918 147704 244924 147756
rect 244976 147704 244982 147756
rect 244936 147620 244964 147704
rect 301498 147676 301504 147688
rect 301459 147648 301504 147676
rect 301498 147636 301504 147648
rect 301556 147636 301562 147688
rect 344094 147636 344100 147688
rect 344152 147676 344158 147688
rect 344278 147676 344284 147688
rect 344152 147648 344284 147676
rect 344152 147636 344158 147648
rect 344278 147636 344284 147648
rect 344336 147636 344342 147688
rect 244366 147568 244372 147620
rect 244424 147568 244430 147620
rect 244918 147568 244924 147620
rect 244976 147568 244982 147620
rect 345290 144916 345296 144968
rect 345348 144956 345354 144968
rect 345382 144956 345388 144968
rect 345348 144928 345388 144956
rect 345348 144916 345354 144928
rect 345382 144916 345388 144928
rect 345440 144916 345446 144968
rect 232038 143596 232044 143608
rect 231999 143568 232044 143596
rect 232038 143556 232044 143568
rect 232096 143556 232102 143608
rect 246390 143596 246396 143608
rect 246351 143568 246396 143596
rect 246390 143556 246396 143568
rect 246448 143556 246454 143608
rect 320910 143556 320916 143608
rect 320968 143596 320974 143608
rect 321094 143596 321100 143608
rect 320968 143568 321100 143596
rect 320968 143556 320974 143568
rect 321094 143556 321100 143568
rect 321152 143556 321158 143608
rect 107470 143528 107476 143540
rect 107431 143500 107476 143528
rect 107470 143488 107476 143500
rect 107528 143488 107534 143540
rect 240686 143528 240692 143540
rect 240647 143500 240692 143528
rect 240686 143488 240692 143500
rect 240744 143488 240750 143540
rect 244366 143488 244372 143540
rect 244424 143528 244430 143540
rect 244458 143528 244464 143540
rect 244424 143500 244464 143528
rect 244424 143488 244430 143500
rect 244458 143488 244464 143500
rect 244516 143488 244522 143540
rect 246022 143528 246028 143540
rect 245983 143500 246028 143528
rect 246022 143488 246028 143500
rect 246080 143488 246086 143540
rect 254670 143488 254676 143540
rect 254728 143528 254734 143540
rect 254854 143528 254860 143540
rect 254728 143500 254860 143528
rect 254728 143488 254734 143500
rect 254854 143488 254860 143500
rect 254912 143488 254918 143540
rect 258810 143528 258816 143540
rect 258771 143500 258816 143528
rect 258810 143488 258816 143500
rect 258868 143488 258874 143540
rect 314286 143488 314292 143540
rect 314344 143488 314350 143540
rect 314378 143488 314384 143540
rect 314436 143528 314442 143540
rect 314436 143500 314481 143528
rect 314436 143488 314442 143500
rect 314194 143420 314200 143472
rect 314252 143420 314258 143472
rect 314212 143336 314240 143420
rect 314304 143404 314332 143488
rect 314286 143352 314292 143404
rect 314344 143352 314350 143404
rect 314194 143284 314200 143336
rect 314252 143284 314258 143336
rect 253017 142239 253075 142245
rect 253017 142205 253029 142239
rect 253063 142236 253075 142239
rect 253198 142236 253204 142248
rect 253063 142208 253204 142236
rect 253063 142205 253075 142208
rect 253017 142199 253075 142205
rect 253198 142196 253204 142208
rect 253256 142196 253262 142248
rect 246390 142168 246396 142180
rect 246351 142140 246396 142168
rect 246390 142128 246396 142140
rect 246448 142128 246454 142180
rect 256970 142128 256976 142180
rect 257028 142168 257034 142180
rect 257338 142168 257344 142180
rect 257028 142140 257344 142168
rect 257028 142128 257034 142140
rect 257338 142128 257344 142140
rect 257396 142128 257402 142180
rect 260282 142128 260288 142180
rect 260340 142128 260346 142180
rect 264514 142168 264520 142180
rect 264475 142140 264520 142168
rect 264514 142128 264520 142140
rect 264572 142128 264578 142180
rect 294690 142128 294696 142180
rect 294748 142168 294754 142180
rect 294782 142168 294788 142180
rect 294748 142140 294788 142168
rect 294748 142128 294754 142140
rect 294782 142128 294788 142140
rect 294840 142128 294846 142180
rect 326154 142128 326160 142180
rect 326212 142168 326218 142180
rect 326338 142168 326344 142180
rect 326212 142140 326344 142168
rect 326212 142128 326218 142140
rect 326338 142128 326344 142140
rect 326396 142128 326402 142180
rect 331766 142168 331772 142180
rect 331727 142140 331772 142168
rect 331766 142128 331772 142140
rect 331824 142128 331830 142180
rect 334526 142168 334532 142180
rect 334487 142140 334532 142168
rect 334526 142128 334532 142140
rect 334584 142128 334590 142180
rect 232038 142100 232044 142112
rect 231999 142072 232044 142100
rect 232038 142060 232044 142072
rect 232096 142060 232102 142112
rect 260300 142044 260328 142128
rect 293310 142100 293316 142112
rect 293271 142072 293316 142100
rect 293310 142060 293316 142072
rect 293368 142060 293374 142112
rect 319622 142100 319628 142112
rect 319583 142072 319628 142100
rect 319622 142060 319628 142072
rect 319680 142060 319686 142112
rect 322290 142060 322296 142112
rect 322348 142060 322354 142112
rect 246390 141992 246396 142044
rect 246448 141992 246454 142044
rect 260282 141992 260288 142044
rect 260340 141992 260346 142044
rect 246408 141905 246436 141992
rect 322308 141976 322336 142060
rect 322290 141924 322296 141976
rect 322348 141924 322354 141976
rect 246393 141899 246451 141905
rect 246393 141865 246405 141899
rect 246439 141865 246451 141899
rect 246393 141859 246451 141865
rect 301866 141080 301872 141092
rect 301827 141052 301872 141080
rect 301866 141040 301872 141052
rect 301924 141040 301930 141092
rect 296073 140811 296131 140817
rect 296073 140777 296085 140811
rect 296119 140808 296131 140811
rect 296162 140808 296168 140820
rect 296119 140780 296168 140808
rect 296119 140777 296131 140780
rect 296073 140771 296131 140777
rect 296162 140768 296168 140780
rect 296220 140768 296226 140820
rect 330386 140768 330392 140820
rect 330444 140808 330450 140820
rect 330481 140811 330539 140817
rect 330481 140808 330493 140811
rect 330444 140780 330493 140808
rect 330444 140768 330450 140780
rect 330481 140777 330493 140780
rect 330527 140777 330539 140811
rect 330481 140771 330539 140777
rect 244918 140740 244924 140752
rect 244879 140712 244924 140740
rect 244918 140700 244924 140712
rect 244976 140700 244982 140752
rect 253198 140740 253204 140752
rect 253159 140712 253204 140740
rect 253198 140700 253204 140712
rect 253256 140700 253262 140752
rect 299014 140740 299020 140752
rect 298975 140712 299020 140740
rect 299014 140700 299020 140712
rect 299072 140700 299078 140752
rect 300302 140740 300308 140752
rect 300263 140712 300308 140740
rect 300302 140700 300308 140712
rect 300360 140700 300366 140752
rect 301498 140700 301504 140752
rect 301556 140740 301562 140752
rect 301774 140740 301780 140752
rect 301556 140712 301780 140740
rect 301556 140700 301562 140712
rect 301774 140700 301780 140712
rect 301832 140700 301838 140752
rect 329006 140740 329012 140752
rect 328967 140712 329012 140740
rect 329006 140700 329012 140712
rect 329064 140700 329070 140752
rect 331766 140740 331772 140752
rect 331727 140712 331772 140740
rect 331766 140700 331772 140712
rect 331824 140700 331830 140752
rect 335814 140700 335820 140752
rect 335872 140740 335878 140752
rect 335909 140743 335967 140749
rect 335909 140740 335921 140743
rect 335872 140712 335921 140740
rect 335872 140700 335878 140712
rect 335909 140709 335921 140712
rect 335955 140709 335967 140743
rect 335909 140703 335967 140709
rect 301866 140672 301872 140684
rect 301827 140644 301872 140672
rect 301866 140632 301872 140644
rect 301924 140632 301930 140684
rect 232406 139340 232412 139392
rect 232464 139380 232470 139392
rect 232590 139380 232596 139392
rect 232464 139352 232596 139380
rect 232464 139340 232470 139352
rect 232590 139340 232596 139352
rect 232648 139340 232654 139392
rect 260190 139380 260196 139392
rect 260151 139352 260196 139380
rect 260190 139340 260196 139352
rect 260248 139340 260254 139392
rect 258813 138635 258871 138641
rect 258813 138601 258825 138635
rect 258859 138632 258871 138635
rect 258902 138632 258908 138644
rect 258859 138604 258908 138632
rect 258859 138601 258871 138604
rect 258813 138595 258871 138601
rect 258902 138592 258908 138604
rect 258960 138592 258966 138644
rect 314378 138496 314384 138508
rect 314339 138468 314384 138496
rect 314378 138456 314384 138468
rect 314436 138456 314442 138508
rect 232590 138048 232596 138100
rect 232648 138088 232654 138100
rect 232682 138088 232688 138100
rect 232648 138060 232688 138088
rect 232648 138048 232654 138060
rect 232682 138048 232688 138060
rect 232740 138048 232746 138100
rect 231210 138020 231216 138032
rect 231171 137992 231216 138020
rect 231210 137980 231216 137992
rect 231268 137980 231274 138032
rect 232406 136552 232412 136604
rect 232464 136552 232470 136604
rect 232424 136465 232452 136552
rect 232409 136459 232467 136465
rect 232409 136425 232421 136459
rect 232455 136425 232467 136459
rect 232409 136419 232467 136425
rect 2774 136348 2780 136400
rect 2832 136388 2838 136400
rect 4798 136388 4804 136400
rect 2832 136360 4804 136388
rect 2832 136348 2838 136360
rect 4798 136348 4804 136360
rect 4856 136348 4862 136400
rect 231210 135368 231216 135380
rect 231171 135340 231216 135368
rect 231210 135328 231216 135340
rect 231268 135328 231274 135380
rect 340138 135300 340144 135312
rect 340064 135272 340144 135300
rect 340064 135244 340092 135272
rect 340138 135260 340144 135272
rect 340196 135260 340202 135312
rect 345290 135260 345296 135312
rect 345348 135300 345354 135312
rect 345382 135300 345388 135312
rect 345348 135272 345388 135300
rect 345348 135260 345354 135272
rect 345382 135260 345388 135272
rect 345440 135260 345446 135312
rect 100662 135192 100668 135244
rect 100720 135232 100726 135244
rect 100846 135232 100852 135244
rect 100720 135204 100852 135232
rect 100720 135192 100726 135204
rect 100846 135192 100852 135204
rect 100904 135192 100910 135244
rect 231210 135192 231216 135244
rect 231268 135232 231274 135244
rect 231394 135232 231400 135244
rect 231268 135204 231400 135232
rect 231268 135192 231274 135204
rect 231394 135192 231400 135204
rect 231452 135192 231458 135244
rect 340046 135192 340052 135244
rect 340104 135192 340110 135244
rect 301774 134552 301780 134564
rect 301735 134524 301780 134552
rect 301774 134512 301780 134524
rect 301832 134512 301838 134564
rect 107470 133940 107476 133952
rect 107431 133912 107476 133940
rect 107470 133900 107476 133912
rect 107528 133900 107534 133952
rect 240686 133940 240692 133952
rect 240647 133912 240692 133940
rect 240686 133900 240692 133912
rect 240744 133900 240750 133952
rect 340046 133872 340052 133884
rect 340007 133844 340052 133872
rect 340046 133832 340052 133844
rect 340104 133832 340110 133884
rect 345382 133832 345388 133884
rect 345440 133872 345446 133884
rect 345566 133872 345572 133884
rect 345440 133844 345572 133872
rect 345440 133832 345446 133844
rect 345566 133832 345572 133844
rect 345624 133832 345630 133884
rect 245838 133288 245844 133340
rect 245896 133328 245902 133340
rect 246025 133331 246083 133337
rect 246025 133328 246037 133331
rect 245896 133300 246037 133328
rect 245896 133288 245902 133300
rect 246025 133297 246037 133300
rect 246071 133297 246083 133331
rect 246025 133291 246083 133297
rect 232041 132515 232099 132521
rect 232041 132481 232053 132515
rect 232087 132512 232099 132515
rect 232130 132512 232136 132524
rect 232087 132484 232136 132512
rect 232087 132481 232099 132484
rect 232041 132475 232099 132481
rect 232130 132472 232136 132484
rect 232188 132472 232194 132524
rect 293310 132512 293316 132524
rect 293271 132484 293316 132512
rect 293310 132472 293316 132484
rect 293368 132472 293374 132524
rect 294782 132472 294788 132524
rect 294840 132512 294846 132524
rect 294874 132512 294880 132524
rect 294840 132484 294880 132512
rect 294840 132472 294846 132484
rect 294874 132472 294880 132484
rect 294932 132472 294938 132524
rect 319622 132512 319628 132524
rect 319583 132484 319628 132512
rect 319622 132472 319628 132484
rect 319680 132472 319686 132524
rect 321002 132472 321008 132524
rect 321060 132512 321066 132524
rect 321094 132512 321100 132524
rect 321060 132484 321100 132512
rect 321060 132472 321066 132484
rect 321094 132472 321100 132484
rect 321152 132472 321158 132524
rect 326154 132472 326160 132524
rect 326212 132512 326218 132524
rect 326246 132512 326252 132524
rect 326212 132484 326252 132512
rect 326212 132472 326218 132484
rect 326246 132472 326252 132484
rect 326304 132472 326310 132524
rect 330386 132472 330392 132524
rect 330444 132512 330450 132524
rect 330478 132512 330484 132524
rect 330444 132484 330484 132512
rect 330444 132472 330450 132484
rect 330478 132472 330484 132484
rect 330536 132472 330542 132524
rect 244921 131223 244979 131229
rect 244921 131189 244933 131223
rect 244967 131220 244979 131223
rect 244967 131192 245148 131220
rect 244967 131189 244979 131192
rect 244921 131183 244979 131189
rect 245120 131164 245148 131192
rect 261478 131180 261484 131232
rect 261536 131220 261542 131232
rect 261570 131220 261576 131232
rect 261536 131192 261576 131220
rect 261536 131180 261542 131192
rect 261570 131180 261576 131192
rect 261628 131180 261634 131232
rect 245102 131112 245108 131164
rect 245160 131112 245166 131164
rect 253198 131152 253204 131164
rect 253159 131124 253204 131152
rect 253198 131112 253204 131124
rect 253256 131112 253262 131164
rect 329009 131155 329067 131161
rect 329009 131121 329021 131155
rect 329055 131152 329067 131155
rect 329190 131152 329196 131164
rect 329055 131124 329196 131152
rect 329055 131121 329067 131124
rect 329009 131115 329067 131121
rect 329190 131112 329196 131124
rect 329248 131112 329254 131164
rect 331766 131152 331772 131164
rect 331727 131124 331772 131152
rect 331766 131112 331772 131124
rect 331824 131112 331830 131164
rect 335906 131112 335912 131164
rect 335964 131152 335970 131164
rect 335964 131124 336009 131152
rect 335964 131112 335970 131124
rect 261478 131084 261484 131096
rect 261439 131056 261484 131084
rect 261478 131044 261484 131056
rect 261536 131044 261542 131096
rect 334437 131087 334495 131093
rect 334437 131053 334449 131087
rect 334483 131084 334495 131087
rect 334526 131084 334532 131096
rect 334483 131056 334532 131084
rect 334483 131053 334495 131056
rect 334437 131047 334495 131053
rect 334526 131044 334532 131056
rect 334584 131044 334590 131096
rect 300302 130744 300308 130756
rect 300263 130716 300308 130744
rect 300302 130704 300308 130716
rect 300360 130704 300366 130756
rect 299014 129860 299020 129872
rect 298975 129832 299020 129860
rect 299014 129820 299020 129832
rect 299072 129820 299078 129872
rect 260193 129795 260251 129801
rect 260193 129761 260205 129795
rect 260239 129792 260251 129795
rect 260282 129792 260288 129804
rect 260239 129764 260288 129792
rect 260239 129761 260251 129764
rect 260193 129755 260251 129761
rect 260282 129752 260288 129764
rect 260340 129752 260346 129804
rect 299014 129724 299020 129736
rect 298975 129696 299020 129724
rect 299014 129684 299020 129696
rect 299072 129684 299078 129736
rect 344094 128324 344100 128376
rect 344152 128364 344158 128376
rect 344278 128364 344284 128376
rect 344152 128336 344284 128364
rect 344152 128324 344158 128336
rect 344278 128324 344284 128336
rect 344336 128324 344342 128376
rect 232866 127072 232872 127084
rect 232700 127044 232872 127072
rect 232700 127016 232728 127044
rect 232866 127032 232872 127044
rect 232924 127032 232930 127084
rect 232682 126964 232688 127016
rect 232740 126964 232746 127016
rect 258810 125604 258816 125656
rect 258868 125644 258874 125656
rect 258902 125644 258908 125656
rect 258868 125616 258908 125644
rect 258868 125604 258874 125616
rect 258902 125604 258908 125616
rect 258960 125604 258966 125656
rect 246390 124216 246396 124228
rect 246351 124188 246396 124216
rect 246390 124176 246396 124188
rect 246448 124176 246454 124228
rect 326246 124176 326252 124228
rect 326304 124216 326310 124228
rect 326338 124216 326344 124228
rect 326304 124188 326344 124216
rect 326304 124176 326310 124188
rect 326338 124176 326344 124188
rect 326396 124176 326402 124228
rect 329098 124176 329104 124228
rect 329156 124216 329162 124228
rect 329190 124216 329196 124228
rect 329156 124188 329196 124216
rect 329156 124176 329162 124188
rect 329190 124176 329196 124188
rect 329248 124176 329254 124228
rect 340049 124219 340107 124225
rect 340049 124185 340061 124219
rect 340095 124216 340107 124219
rect 340138 124216 340144 124228
rect 340095 124188 340144 124216
rect 340095 124185 340107 124188
rect 340049 124179 340107 124185
rect 340138 124176 340144 124188
rect 340196 124176 340202 124228
rect 107470 124148 107476 124160
rect 107431 124120 107476 124148
rect 107470 124108 107476 124120
rect 107528 124108 107534 124160
rect 317138 124148 317144 124160
rect 317099 124120 317144 124148
rect 317138 124108 317144 124120
rect 317196 124108 317202 124160
rect 317322 124148 317328 124160
rect 317283 124120 317328 124148
rect 317322 124108 317328 124120
rect 317380 124108 317386 124160
rect 345290 124108 345296 124160
rect 345348 124108 345354 124160
rect 577498 124108 577504 124160
rect 577556 124148 577562 124160
rect 579614 124148 579620 124160
rect 577556 124120 579620 124148
rect 577556 124108 577562 124120
rect 579614 124108 579620 124120
rect 579672 124108 579678 124160
rect 314378 124040 314384 124092
rect 314436 124040 314442 124092
rect 345308 124080 345336 124108
rect 345382 124080 345388 124092
rect 345308 124052 345388 124080
rect 345382 124040 345388 124052
rect 345440 124040 345446 124092
rect 314396 123956 314424 124040
rect 314378 123904 314384 123956
rect 314436 123904 314442 123956
rect 321094 122924 321100 122936
rect 320928 122896 321100 122924
rect 320928 122868 320956 122896
rect 321094 122884 321100 122896
rect 321152 122884 321158 122936
rect 322290 122924 322296 122936
rect 322216 122896 322296 122924
rect 294690 122816 294696 122868
rect 294748 122856 294754 122868
rect 294782 122856 294788 122868
rect 294748 122828 294788 122856
rect 294748 122816 294754 122828
rect 294782 122816 294788 122828
rect 294840 122816 294846 122868
rect 320910 122816 320916 122868
rect 320968 122816 320974 122868
rect 244366 122788 244372 122800
rect 244327 122760 244372 122788
rect 244366 122748 244372 122760
rect 244424 122748 244430 122800
rect 253014 122748 253020 122800
rect 253072 122788 253078 122800
rect 253109 122791 253167 122797
rect 253109 122788 253121 122791
rect 253072 122760 253121 122788
rect 253072 122748 253078 122760
rect 253109 122757 253121 122760
rect 253155 122757 253167 122791
rect 253109 122751 253167 122757
rect 254673 122791 254731 122797
rect 254673 122757 254685 122791
rect 254719 122788 254731 122791
rect 254762 122788 254768 122800
rect 254719 122760 254768 122788
rect 254719 122757 254731 122760
rect 254673 122751 254731 122757
rect 254762 122748 254768 122760
rect 254820 122748 254826 122800
rect 257154 122788 257160 122800
rect 257115 122760 257160 122788
rect 257154 122748 257160 122760
rect 257212 122748 257218 122800
rect 264514 122748 264520 122800
rect 264572 122788 264578 122800
rect 264609 122791 264667 122797
rect 264609 122788 264621 122791
rect 264572 122760 264621 122788
rect 264572 122748 264578 122760
rect 264609 122757 264621 122760
rect 264655 122757 264667 122791
rect 265802 122788 265808 122800
rect 265763 122760 265808 122788
rect 264609 122751 264667 122757
rect 265802 122748 265808 122760
rect 265860 122748 265866 122800
rect 319622 122748 319628 122800
rect 319680 122748 319686 122800
rect 261478 122720 261484 122732
rect 261439 122692 261484 122720
rect 261478 122680 261484 122692
rect 261536 122680 261542 122732
rect 319640 122661 319668 122748
rect 322216 122720 322244 122896
rect 322290 122884 322296 122896
rect 322348 122884 322354 122936
rect 335722 122884 335728 122936
rect 335780 122924 335786 122936
rect 335906 122924 335912 122936
rect 335780 122896 335912 122924
rect 335780 122884 335786 122896
rect 335906 122884 335912 122896
rect 335964 122884 335970 122936
rect 335722 122748 335728 122800
rect 335780 122788 335786 122800
rect 335814 122788 335820 122800
rect 335780 122760 335820 122788
rect 335780 122748 335786 122760
rect 335814 122748 335820 122760
rect 335872 122748 335878 122800
rect 322382 122720 322388 122732
rect 322216 122692 322388 122720
rect 322382 122680 322388 122692
rect 322440 122680 322446 122732
rect 319625 122655 319683 122661
rect 319625 122621 319637 122655
rect 319671 122621 319683 122655
rect 319625 122615 319683 122621
rect 301774 121496 301780 121508
rect 301735 121468 301780 121496
rect 301774 121456 301780 121468
rect 301832 121456 301838 121508
rect 334437 121499 334495 121505
rect 334437 121465 334449 121499
rect 334483 121496 334495 121499
rect 334526 121496 334532 121508
rect 334483 121468 334532 121496
rect 334483 121465 334495 121468
rect 334437 121459 334495 121465
rect 334526 121456 334532 121468
rect 334584 121456 334590 121508
rect 245013 121431 245071 121437
rect 245013 121397 245025 121431
rect 245059 121428 245071 121431
rect 245102 121428 245108 121440
rect 245059 121400 245108 121428
rect 245059 121397 245071 121400
rect 245013 121391 245071 121397
rect 245102 121388 245108 121400
rect 245160 121388 245166 121440
rect 261478 121388 261484 121440
rect 261536 121388 261542 121440
rect 331766 121428 331772 121440
rect 331727 121400 331772 121428
rect 331766 121388 331772 121400
rect 331824 121388 331830 121440
rect 261496 121301 261524 121388
rect 261481 121295 261539 121301
rect 261481 121261 261493 121295
rect 261527 121261 261539 121295
rect 261481 121255 261539 121261
rect 299014 120204 299020 120216
rect 298975 120176 299020 120204
rect 299014 120164 299020 120176
rect 299072 120164 299078 120216
rect 298925 120071 298983 120077
rect 298925 120037 298937 120071
rect 298971 120068 298983 120071
rect 299014 120068 299020 120080
rect 298971 120040 299020 120068
rect 298971 120037 298983 120040
rect 298925 120031 298983 120037
rect 299014 120028 299020 120040
rect 299072 120028 299078 120080
rect 300213 120071 300271 120077
rect 300213 120037 300225 120071
rect 300259 120068 300271 120071
rect 300302 120068 300308 120080
rect 300259 120040 300308 120068
rect 300259 120037 300271 120040
rect 300213 120031 300271 120037
rect 300302 120028 300308 120040
rect 300360 120028 300366 120080
rect 301685 120071 301743 120077
rect 301685 120037 301697 120071
rect 301731 120068 301743 120071
rect 301774 120068 301780 120080
rect 301731 120040 301780 120068
rect 301731 120037 301743 120040
rect 301685 120031 301743 120037
rect 301774 120028 301780 120040
rect 301832 120028 301838 120080
rect 231210 118708 231216 118720
rect 231171 118680 231216 118708
rect 231210 118668 231216 118680
rect 231268 118668 231274 118720
rect 232406 118708 232412 118720
rect 232367 118680 232412 118708
rect 232406 118668 232412 118680
rect 232464 118668 232470 118720
rect 232590 118668 232596 118720
rect 232648 118708 232654 118720
rect 232682 118708 232688 118720
rect 232648 118680 232688 118708
rect 232648 118668 232654 118680
rect 232682 118668 232688 118680
rect 232740 118668 232746 118720
rect 263042 118028 263048 118040
rect 263003 118000 263048 118028
rect 263042 117988 263048 118000
rect 263100 117988 263106 118040
rect 317138 117552 317144 117564
rect 317099 117524 317144 117552
rect 317138 117512 317144 117524
rect 317196 117512 317202 117564
rect 232682 117240 232688 117292
rect 232740 117240 232746 117292
rect 232700 117212 232728 117240
rect 232866 117212 232872 117224
rect 232700 117184 232872 117212
rect 232866 117172 232872 117184
rect 232924 117172 232930 117224
rect 231210 116056 231216 116068
rect 231171 116028 231216 116056
rect 231210 116016 231216 116028
rect 231268 116016 231274 116068
rect 100662 115920 100668 115932
rect 100623 115892 100668 115920
rect 100662 115880 100668 115892
rect 100720 115880 100726 115932
rect 231210 115920 231216 115932
rect 231171 115892 231216 115920
rect 231210 115880 231216 115892
rect 231268 115880 231274 115932
rect 258902 115920 258908 115932
rect 258863 115892 258908 115920
rect 258902 115880 258908 115892
rect 258960 115880 258966 115932
rect 260374 115920 260380 115932
rect 260335 115892 260380 115920
rect 260374 115880 260380 115892
rect 260432 115880 260438 115932
rect 317322 115580 317328 115592
rect 317283 115552 317328 115580
rect 317322 115540 317328 115552
rect 317380 115540 317386 115592
rect 339957 115515 340015 115521
rect 339957 115481 339969 115515
rect 340003 115512 340015 115515
rect 340138 115512 340144 115524
rect 340003 115484 340144 115512
rect 340003 115481 340015 115484
rect 339957 115475 340015 115481
rect 340138 115472 340144 115484
rect 340196 115472 340202 115524
rect 107470 114560 107476 114572
rect 107431 114532 107476 114560
rect 107470 114520 107476 114532
rect 107528 114520 107534 114572
rect 329006 114520 329012 114572
rect 329064 114560 329070 114572
rect 329098 114560 329104 114572
rect 329064 114532 329104 114560
rect 329064 114520 329070 114532
rect 329098 114520 329104 114532
rect 329156 114520 329162 114572
rect 316954 114492 316960 114504
rect 316915 114464 316960 114492
rect 316954 114452 316960 114464
rect 317012 114452 317018 114504
rect 317138 114492 317144 114504
rect 317099 114464 317144 114492
rect 317138 114452 317144 114464
rect 317196 114452 317202 114504
rect 317322 114492 317328 114504
rect 317283 114464 317328 114492
rect 317322 114452 317328 114464
rect 317380 114452 317386 114504
rect 326154 114452 326160 114504
rect 326212 114492 326218 114504
rect 326338 114492 326344 114504
rect 326212 114464 326344 114492
rect 326212 114452 326218 114464
rect 326338 114452 326344 114464
rect 326396 114452 326402 114504
rect 317230 114424 317236 114436
rect 317191 114396 317236 114424
rect 317230 114384 317236 114396
rect 317288 114384 317294 114436
rect 244369 113203 244427 113209
rect 244369 113169 244381 113203
rect 244415 113200 244427 113203
rect 244458 113200 244464 113212
rect 244415 113172 244464 113200
rect 244415 113169 244427 113172
rect 244369 113163 244427 113169
rect 244458 113160 244464 113172
rect 244516 113160 244522 113212
rect 257154 113160 257160 113212
rect 257212 113200 257218 113212
rect 257212 113172 257257 113200
rect 257212 113160 257218 113172
rect 264514 113160 264520 113212
rect 264572 113200 264578 113212
rect 264609 113203 264667 113209
rect 264609 113200 264621 113203
rect 264572 113172 264621 113200
rect 264572 113160 264578 113172
rect 264609 113169 264621 113172
rect 264655 113169 264667 113203
rect 265802 113200 265808 113212
rect 265763 113172 265808 113200
rect 264609 113163 264667 113169
rect 265802 113160 265808 113172
rect 265860 113160 265866 113212
rect 319622 113200 319628 113212
rect 319583 113172 319628 113200
rect 319622 113160 319628 113172
rect 319680 113160 319686 113212
rect 245013 113135 245071 113141
rect 245013 113101 245025 113135
rect 245059 113132 245071 113135
rect 245102 113132 245108 113144
rect 245059 113104 245108 113132
rect 245059 113101 245071 113104
rect 245013 113095 245071 113101
rect 245102 113092 245108 113104
rect 245160 113092 245166 113144
rect 294782 113132 294788 113144
rect 294743 113104 294788 113132
rect 294782 113092 294788 113104
rect 294840 113092 294846 113144
rect 326154 113132 326160 113144
rect 326115 113104 326160 113132
rect 326154 113092 326160 113104
rect 326212 113092 326218 113144
rect 335814 113132 335820 113144
rect 335775 113104 335820 113132
rect 335814 113092 335820 113104
rect 335872 113092 335878 113144
rect 244369 113067 244427 113073
rect 244369 113033 244381 113067
rect 244415 113064 244427 113067
rect 244458 113064 244464 113076
rect 244415 113036 244464 113064
rect 244415 113033 244427 113036
rect 244369 113027 244427 113033
rect 244458 113024 244464 113036
rect 244516 113024 244522 113076
rect 261478 111840 261484 111852
rect 261439 111812 261484 111840
rect 261478 111800 261484 111812
rect 261536 111800 261542 111852
rect 331766 111840 331772 111852
rect 331727 111812 331772 111840
rect 331766 111800 331772 111812
rect 331824 111800 331830 111852
rect 232038 111732 232044 111784
rect 232096 111772 232102 111784
rect 232130 111772 232136 111784
rect 232096 111744 232136 111772
rect 232096 111732 232102 111744
rect 232130 111732 232136 111744
rect 232188 111732 232194 111784
rect 334526 111772 334532 111784
rect 334487 111744 334532 111772
rect 334526 111732 334532 111744
rect 334584 111732 334590 111784
rect 317322 109732 317328 109744
rect 317283 109704 317328 109732
rect 317322 109692 317328 109704
rect 317380 109692 317386 109744
rect 344094 109012 344100 109064
rect 344152 109052 344158 109064
rect 344278 109052 344284 109064
rect 344152 109024 344284 109052
rect 344152 109012 344158 109024
rect 344278 109012 344284 109024
rect 344336 109012 344342 109064
rect 3326 108944 3332 108996
rect 3384 108984 3390 108996
rect 31018 108984 31024 108996
rect 3384 108956 31024 108984
rect 3384 108944 3390 108956
rect 31018 108944 31024 108956
rect 31076 108944 31082 108996
rect 339957 108987 340015 108993
rect 339957 108953 339969 108987
rect 340003 108984 340015 108987
rect 340046 108984 340052 108996
rect 340003 108956 340052 108984
rect 340003 108953 340015 108956
rect 339957 108947 340015 108953
rect 340046 108944 340052 108956
rect 340104 108944 340110 108996
rect 253109 108375 253167 108381
rect 253109 108341 253121 108375
rect 253155 108372 253167 108375
rect 253198 108372 253204 108384
rect 253155 108344 253204 108372
rect 253155 108341 253167 108344
rect 253109 108335 253167 108341
rect 253198 108332 253204 108344
rect 253256 108332 253262 108384
rect 317138 107624 317144 107636
rect 317099 107596 317144 107624
rect 317138 107584 317144 107596
rect 317196 107584 317202 107636
rect 232314 107012 232320 107024
rect 232275 106984 232320 107012
rect 232314 106972 232320 106984
rect 232372 106972 232378 107024
rect 244918 106972 244924 107024
rect 244976 107012 244982 107024
rect 245102 107012 245108 107024
rect 244976 106984 245108 107012
rect 244976 106972 244982 106984
rect 245102 106972 245108 106984
rect 245160 106972 245166 107024
rect 297453 106947 297511 106953
rect 297453 106913 297465 106947
rect 297499 106944 297511 106947
rect 297542 106944 297548 106956
rect 297499 106916 297548 106944
rect 297499 106913 297511 106916
rect 297453 106907 297511 106913
rect 297542 106904 297548 106916
rect 297600 106904 297606 106956
rect 100662 106332 100668 106344
rect 100623 106304 100668 106332
rect 100662 106292 100668 106304
rect 100720 106292 100726 106344
rect 231210 106332 231216 106344
rect 231171 106304 231216 106332
rect 231210 106292 231216 106304
rect 231268 106292 231274 106344
rect 258902 106332 258908 106344
rect 258863 106304 258908 106332
rect 258902 106292 258908 106304
rect 258960 106292 258966 106344
rect 260374 106332 260380 106344
rect 260335 106304 260380 106332
rect 260374 106292 260380 106304
rect 260432 106292 260438 106344
rect 317230 106128 317236 106140
rect 317191 106100 317236 106128
rect 317230 106088 317236 106100
rect 317288 106088 317294 106140
rect 321094 106060 321100 106072
rect 321055 106032 321100 106060
rect 321094 106020 321100 106032
rect 321152 106020 321158 106072
rect 246482 104864 246488 104916
rect 246540 104904 246546 104916
rect 246574 104904 246580 104916
rect 246540 104876 246580 104904
rect 246540 104864 246546 104876
rect 246574 104864 246580 104876
rect 246632 104864 246638 104916
rect 254670 104904 254676 104916
rect 254631 104876 254676 104904
rect 254670 104864 254676 104876
rect 254728 104864 254734 104916
rect 263042 104904 263048 104916
rect 263003 104876 263048 104904
rect 263042 104864 263048 104876
rect 263100 104864 263106 104916
rect 316954 104904 316960 104916
rect 316915 104876 316960 104904
rect 316954 104864 316960 104876
rect 317012 104864 317018 104916
rect 322290 104864 322296 104916
rect 322348 104904 322354 104916
rect 322382 104904 322388 104916
rect 322348 104876 322388 104904
rect 322348 104864 322354 104876
rect 322382 104864 322388 104876
rect 322440 104864 322446 104916
rect 107470 104836 107476 104848
rect 107431 104808 107476 104836
rect 107470 104796 107476 104808
rect 107528 104796 107534 104848
rect 244366 103612 244372 103624
rect 244327 103584 244372 103612
rect 244366 103572 244372 103584
rect 244424 103572 244430 103624
rect 261478 103612 261484 103624
rect 261404 103584 261484 103612
rect 261404 103556 261432 103584
rect 261478 103572 261484 103584
rect 261536 103572 261542 103624
rect 321186 103612 321192 103624
rect 321112 103584 321192 103612
rect 261386 103504 261392 103556
rect 261444 103504 261450 103556
rect 294782 103544 294788 103556
rect 294743 103516 294788 103544
rect 294782 103504 294788 103516
rect 294840 103504 294846 103556
rect 295978 103504 295984 103556
rect 296036 103544 296042 103556
rect 296070 103544 296076 103556
rect 296036 103516 296076 103544
rect 296036 103504 296042 103516
rect 296070 103504 296076 103516
rect 296128 103504 296134 103556
rect 321112 103488 321140 103584
rect 321186 103572 321192 103584
rect 321244 103572 321250 103624
rect 329006 103612 329012 103624
rect 328932 103584 329012 103612
rect 328932 103556 328960 103584
rect 329006 103572 329012 103584
rect 329064 103572 329070 103624
rect 330478 103612 330484 103624
rect 330404 103584 330484 103612
rect 330404 103556 330432 103584
rect 330478 103572 330484 103584
rect 330536 103572 330542 103624
rect 335814 103612 335820 103624
rect 335775 103584 335820 103612
rect 335814 103572 335820 103584
rect 335872 103572 335878 103624
rect 326157 103547 326215 103553
rect 326157 103513 326169 103547
rect 326203 103544 326215 103547
rect 326246 103544 326252 103556
rect 326203 103516 326252 103544
rect 326203 103513 326215 103516
rect 326157 103507 326215 103513
rect 326246 103504 326252 103516
rect 326304 103504 326310 103556
rect 328914 103504 328920 103556
rect 328972 103504 328978 103556
rect 330386 103504 330392 103556
rect 330444 103504 330450 103556
rect 244366 103436 244372 103488
rect 244424 103476 244430 103488
rect 244642 103476 244648 103488
rect 244424 103448 244648 103476
rect 244424 103436 244430 103448
rect 244642 103436 244648 103448
rect 244700 103436 244706 103488
rect 253198 103476 253204 103488
rect 253159 103448 253204 103476
rect 253198 103436 253204 103448
rect 253256 103436 253262 103488
rect 258902 103476 258908 103488
rect 258863 103448 258908 103476
rect 258902 103436 258908 103448
rect 258960 103436 258966 103488
rect 263042 103476 263048 103488
rect 263003 103448 263048 103476
rect 263042 103436 263048 103448
rect 263100 103436 263106 103488
rect 264425 103479 264483 103485
rect 264425 103445 264437 103479
rect 264471 103476 264483 103479
rect 264514 103476 264520 103488
rect 264471 103448 264520 103476
rect 264471 103445 264483 103448
rect 264425 103439 264483 103445
rect 264514 103436 264520 103448
rect 264572 103436 264578 103488
rect 265713 103479 265771 103485
rect 265713 103445 265725 103479
rect 265759 103476 265771 103479
rect 265802 103476 265808 103488
rect 265759 103448 265808 103476
rect 265759 103445 265771 103448
rect 265713 103439 265771 103445
rect 265802 103436 265808 103448
rect 265860 103436 265866 103488
rect 293310 103476 293316 103488
rect 293271 103448 293316 103476
rect 293310 103436 293316 103448
rect 293368 103436 293374 103488
rect 319622 103476 319628 103488
rect 319583 103448 319628 103476
rect 319622 103436 319628 103448
rect 319680 103436 319686 103488
rect 321094 103436 321100 103488
rect 321152 103436 321158 103488
rect 321278 103436 321284 103488
rect 321336 103436 321342 103488
rect 322290 103476 322296 103488
rect 322251 103448 322296 103476
rect 322290 103436 322296 103448
rect 322348 103436 322354 103488
rect 331766 103436 331772 103488
rect 331824 103476 331830 103488
rect 331858 103476 331864 103488
rect 331824 103448 331864 103476
rect 331824 103436 331830 103448
rect 331858 103436 331864 103448
rect 331916 103436 331922 103488
rect 333238 103436 333244 103488
rect 333296 103476 333302 103488
rect 333330 103476 333336 103488
rect 333296 103448 333336 103476
rect 333296 103436 333302 103448
rect 333330 103436 333336 103448
rect 333388 103436 333394 103488
rect 335814 103436 335820 103488
rect 335872 103476 335878 103488
rect 335909 103479 335967 103485
rect 335909 103476 335921 103479
rect 335872 103448 335921 103476
rect 335872 103436 335878 103448
rect 335909 103445 335921 103448
rect 335955 103445 335967 103479
rect 335909 103439 335967 103445
rect 321296 103284 321324 103436
rect 321278 103232 321284 103284
rect 321336 103232 321342 103284
rect 334526 102252 334532 102264
rect 334487 102224 334532 102252
rect 334526 102212 334532 102224
rect 334584 102212 334590 102264
rect 298922 102184 298928 102196
rect 298883 102156 298928 102184
rect 298922 102144 298928 102156
rect 298980 102144 298986 102196
rect 300210 102184 300216 102196
rect 300171 102156 300216 102184
rect 300210 102144 300216 102156
rect 300268 102144 300274 102196
rect 301682 102184 301688 102196
rect 301643 102156 301688 102184
rect 301682 102144 301688 102156
rect 301740 102144 301746 102196
rect 232130 102116 232136 102128
rect 232091 102088 232136 102116
rect 232130 102076 232136 102088
rect 232188 102076 232194 102128
rect 328914 102116 328920 102128
rect 328875 102088 328920 102116
rect 328914 102076 328920 102088
rect 328972 102076 328978 102128
rect 334526 102116 334532 102128
rect 334487 102088 334532 102116
rect 334526 102076 334532 102088
rect 334584 102076 334590 102128
rect 297450 100756 297456 100768
rect 297411 100728 297456 100756
rect 297450 100716 297456 100728
rect 297508 100716 297514 100768
rect 261386 99764 261392 99816
rect 261444 99804 261450 99816
rect 261573 99807 261631 99813
rect 261573 99804 261585 99807
rect 261444 99776 261585 99804
rect 261444 99764 261450 99776
rect 261573 99773 261585 99776
rect 261619 99773 261631 99807
rect 261573 99767 261631 99773
rect 232682 99424 232688 99476
rect 232740 99424 232746 99476
rect 246301 99467 246359 99473
rect 246301 99433 246313 99467
rect 246347 99464 246359 99467
rect 246482 99464 246488 99476
rect 246347 99436 246488 99464
rect 246347 99433 246359 99436
rect 246301 99427 246359 99433
rect 246482 99424 246488 99436
rect 246540 99424 246546 99476
rect 231210 99396 231216 99408
rect 231171 99368 231216 99396
rect 231210 99356 231216 99368
rect 231268 99356 231274 99408
rect 232700 99340 232728 99424
rect 244918 99356 244924 99408
rect 244976 99396 244982 99408
rect 244976 99368 245056 99396
rect 244976 99356 244982 99368
rect 245028 99340 245056 99368
rect 232682 99288 232688 99340
rect 232740 99288 232746 99340
rect 245010 99288 245016 99340
rect 245068 99288 245074 99340
rect 231210 96744 231216 96756
rect 231171 96716 231216 96744
rect 231210 96704 231216 96716
rect 231268 96704 231274 96756
rect 297450 96636 297456 96688
rect 297508 96636 297514 96688
rect 345290 96636 345296 96688
rect 345348 96676 345354 96688
rect 345382 96676 345388 96688
rect 345348 96648 345388 96676
rect 345348 96636 345354 96648
rect 345382 96636 345388 96648
rect 345440 96636 345446 96688
rect 100662 96608 100668 96620
rect 100623 96580 100668 96608
rect 100662 96568 100668 96580
rect 100720 96568 100726 96620
rect 297468 96540 297496 96636
rect 297542 96540 297548 96552
rect 297468 96512 297548 96540
rect 297542 96500 297548 96512
rect 297600 96500 297606 96552
rect 294782 95316 294788 95328
rect 294708 95288 294788 95316
rect 107470 95248 107476 95260
rect 107431 95220 107476 95248
rect 107470 95208 107476 95220
rect 107528 95208 107534 95260
rect 254670 95208 254676 95260
rect 254728 95248 254734 95260
rect 254762 95248 254768 95260
rect 254728 95220 254768 95248
rect 254728 95208 254734 95220
rect 254762 95208 254768 95220
rect 254820 95208 254826 95260
rect 294708 95192 294736 95288
rect 294782 95276 294788 95288
rect 294840 95276 294846 95328
rect 246298 95180 246304 95192
rect 246259 95152 246304 95180
rect 246298 95140 246304 95152
rect 246356 95140 246362 95192
rect 253198 95180 253204 95192
rect 253159 95152 253204 95180
rect 253198 95140 253204 95152
rect 253256 95140 253262 95192
rect 257065 95183 257123 95189
rect 257065 95149 257077 95183
rect 257111 95180 257123 95183
rect 257154 95180 257160 95192
rect 257111 95152 257160 95180
rect 257111 95149 257123 95152
rect 257065 95143 257123 95149
rect 257154 95140 257160 95152
rect 257212 95140 257218 95192
rect 265710 95180 265716 95192
rect 265671 95152 265716 95180
rect 265710 95140 265716 95152
rect 265768 95140 265774 95192
rect 294690 95140 294696 95192
rect 294748 95140 294754 95192
rect 340046 95180 340052 95192
rect 340007 95152 340052 95180
rect 340046 95140 340052 95152
rect 340104 95140 340110 95192
rect 232314 93888 232320 93900
rect 232275 93860 232320 93888
rect 232314 93848 232320 93860
rect 232372 93848 232378 93900
rect 258902 93888 258908 93900
rect 258863 93860 258908 93888
rect 258902 93848 258908 93860
rect 258960 93848 258966 93900
rect 263042 93888 263048 93900
rect 263003 93860 263048 93888
rect 263042 93848 263048 93860
rect 263100 93848 263106 93900
rect 264422 93888 264428 93900
rect 264383 93860 264428 93888
rect 264422 93848 264428 93860
rect 264480 93848 264486 93900
rect 293310 93888 293316 93900
rect 293271 93860 293316 93888
rect 293310 93848 293316 93860
rect 293368 93848 293374 93900
rect 295978 93848 295984 93900
rect 296036 93888 296042 93900
rect 296070 93888 296076 93900
rect 296036 93860 296076 93888
rect 296036 93848 296042 93860
rect 296070 93848 296076 93860
rect 296128 93848 296134 93900
rect 319622 93888 319628 93900
rect 319583 93860 319628 93888
rect 319622 93848 319628 93860
rect 319680 93848 319686 93900
rect 321094 93888 321100 93900
rect 321055 93860 321100 93888
rect 321094 93848 321100 93860
rect 321152 93848 321158 93900
rect 322293 93891 322351 93897
rect 322293 93857 322305 93891
rect 322339 93888 322351 93891
rect 322382 93888 322388 93900
rect 322339 93860 322388 93888
rect 322339 93857 322351 93860
rect 322293 93851 322351 93857
rect 322382 93848 322388 93860
rect 322440 93848 322446 93900
rect 330386 93848 330392 93900
rect 330444 93888 330450 93900
rect 330478 93888 330484 93900
rect 330444 93860 330484 93888
rect 330444 93848 330450 93860
rect 330478 93848 330484 93860
rect 330536 93848 330542 93900
rect 335906 93848 335912 93900
rect 335964 93888 335970 93900
rect 335964 93860 336009 93888
rect 335964 93848 335970 93860
rect 298922 93780 298928 93832
rect 298980 93780 298986 93832
rect 300210 93780 300216 93832
rect 300268 93780 300274 93832
rect 301682 93780 301688 93832
rect 301740 93780 301746 93832
rect 298940 93752 298968 93780
rect 299014 93752 299020 93764
rect 298940 93724 299020 93752
rect 299014 93712 299020 93724
rect 299072 93712 299078 93764
rect 300228 93752 300256 93780
rect 300302 93752 300308 93764
rect 300228 93724 300308 93752
rect 300302 93712 300308 93724
rect 300360 93712 300366 93764
rect 301700 93752 301728 93780
rect 301774 93752 301780 93764
rect 301700 93724 301780 93752
rect 301774 93712 301780 93724
rect 301832 93712 301838 93764
rect 232130 92528 232136 92540
rect 232091 92500 232136 92528
rect 232130 92488 232136 92500
rect 232188 92488 232194 92540
rect 328917 92531 328975 92537
rect 328917 92497 328929 92531
rect 328963 92528 328975 92531
rect 329190 92528 329196 92540
rect 328963 92500 329196 92528
rect 328963 92497 328975 92500
rect 328917 92491 328975 92497
rect 329190 92488 329196 92500
rect 329248 92488 329254 92540
rect 334529 92531 334587 92537
rect 334529 92497 334541 92531
rect 334575 92528 334587 92531
rect 334618 92528 334624 92540
rect 334575 92500 334624 92528
rect 334575 92497 334587 92500
rect 334529 92491 334587 92497
rect 334618 92488 334624 92500
rect 334676 92488 334682 92540
rect 263042 89768 263048 89820
rect 263100 89768 263106 89820
rect 232314 89740 232320 89752
rect 232275 89712 232320 89740
rect 232314 89700 232320 89712
rect 232372 89700 232378 89752
rect 263060 89684 263088 89768
rect 344094 89700 344100 89752
rect 344152 89740 344158 89752
rect 344278 89740 344284 89752
rect 344152 89712 344284 89740
rect 344152 89700 344158 89712
rect 344278 89700 344284 89712
rect 344336 89700 344342 89752
rect 263042 89632 263048 89684
rect 263100 89632 263106 89684
rect 296622 89060 296628 89072
rect 296583 89032 296628 89060
rect 296622 89020 296628 89032
rect 296680 89020 296686 89072
rect 379422 87116 379428 87168
rect 379480 87156 379486 87168
rect 386322 87156 386328 87168
rect 379480 87128 386328 87156
rect 379480 87116 379486 87128
rect 386322 87116 386328 87128
rect 386380 87116 386386 87168
rect 100662 87020 100668 87032
rect 100623 86992 100668 87020
rect 100662 86980 100668 86992
rect 100720 86980 100726 87032
rect 246022 86980 246028 87032
rect 246080 86980 246086 87032
rect 246040 86884 246068 86980
rect 249702 86912 249708 86964
rect 249760 86952 249766 86964
rect 252094 86952 252100 86964
rect 249760 86924 252100 86952
rect 249760 86912 249766 86924
rect 252094 86912 252100 86924
rect 252152 86912 252158 86964
rect 246114 86884 246120 86896
rect 246040 86856 246120 86884
rect 246114 86844 246120 86856
rect 246172 86844 246178 86896
rect 296622 86884 296628 86896
rect 296583 86856 296628 86884
rect 296622 86844 296628 86856
rect 296680 86844 296686 86896
rect 253017 85663 253075 85669
rect 253017 85629 253029 85663
rect 253063 85660 253075 85663
rect 253198 85660 253204 85672
rect 253063 85632 253204 85660
rect 253063 85629 253075 85632
rect 253017 85623 253075 85629
rect 253198 85620 253204 85632
rect 253256 85620 253262 85672
rect 244458 85552 244464 85604
rect 244516 85592 244522 85604
rect 244642 85592 244648 85604
rect 244516 85564 244648 85592
rect 244516 85552 244522 85564
rect 244642 85552 244648 85564
rect 244700 85552 244706 85604
rect 246298 85552 246304 85604
rect 246356 85592 246362 85604
rect 246390 85592 246396 85604
rect 246356 85564 246396 85592
rect 246356 85552 246362 85564
rect 246390 85552 246396 85564
rect 246448 85552 246454 85604
rect 257062 85592 257068 85604
rect 257023 85564 257068 85592
rect 257062 85552 257068 85564
rect 257120 85552 257126 85604
rect 260282 85552 260288 85604
rect 260340 85592 260346 85604
rect 260374 85592 260380 85604
rect 260340 85564 260380 85592
rect 260340 85552 260346 85564
rect 260374 85552 260380 85564
rect 260432 85552 260438 85604
rect 264422 85552 264428 85604
rect 264480 85592 264486 85604
rect 264514 85592 264520 85604
rect 264480 85564 264520 85592
rect 264480 85552 264486 85564
rect 264514 85552 264520 85564
rect 264572 85552 264578 85604
rect 265710 85552 265716 85604
rect 265768 85592 265774 85604
rect 265802 85592 265808 85604
rect 265768 85564 265808 85592
rect 265768 85552 265774 85564
rect 265802 85552 265808 85564
rect 265860 85552 265866 85604
rect 294690 85552 294696 85604
rect 294748 85592 294754 85604
rect 294782 85592 294788 85604
rect 294748 85564 294788 85592
rect 294748 85552 294754 85564
rect 294782 85552 294788 85564
rect 294840 85552 294846 85604
rect 322290 85552 322296 85604
rect 322348 85592 322354 85604
rect 322382 85592 322388 85604
rect 322348 85564 322388 85592
rect 322348 85552 322354 85564
rect 322382 85552 322388 85564
rect 322440 85552 322446 85604
rect 331766 85552 331772 85604
rect 331824 85592 331830 85604
rect 331858 85592 331864 85604
rect 331824 85564 331864 85592
rect 331824 85552 331830 85564
rect 331858 85552 331864 85564
rect 331916 85552 331922 85604
rect 333238 85552 333244 85604
rect 333296 85592 333302 85604
rect 333330 85592 333336 85604
rect 333296 85564 333336 85592
rect 333296 85552 333302 85564
rect 333330 85552 333336 85564
rect 333388 85552 333394 85604
rect 340049 85595 340107 85601
rect 340049 85561 340061 85595
rect 340095 85592 340107 85595
rect 340138 85592 340144 85604
rect 340095 85564 340144 85592
rect 340095 85561 340107 85564
rect 340049 85555 340107 85561
rect 340138 85552 340144 85564
rect 340196 85552 340202 85604
rect 107470 85524 107476 85536
rect 107431 85496 107476 85524
rect 107470 85484 107476 85496
rect 107528 85484 107534 85536
rect 261573 85527 261631 85533
rect 261573 85493 261585 85527
rect 261619 85524 261631 85527
rect 261662 85524 261668 85536
rect 261619 85496 261668 85524
rect 261619 85493 261631 85496
rect 261573 85487 261631 85493
rect 261662 85484 261668 85496
rect 261720 85484 261726 85536
rect 232222 85348 232228 85400
rect 232280 85348 232286 85400
rect 232240 85264 232268 85348
rect 232222 85212 232228 85264
rect 232280 85212 232286 85264
rect 320821 84303 320879 84309
rect 320821 84269 320833 84303
rect 320867 84300 320879 84303
rect 321094 84300 321100 84312
rect 320867 84272 321100 84300
rect 320867 84269 320879 84272
rect 320821 84263 320879 84269
rect 321094 84260 321100 84272
rect 321152 84260 321158 84312
rect 253014 84232 253020 84244
rect 252975 84204 253020 84232
rect 253014 84192 253020 84204
rect 253072 84192 253078 84244
rect 258718 84192 258724 84244
rect 258776 84232 258782 84244
rect 258902 84232 258908 84244
rect 258776 84204 258908 84232
rect 258776 84192 258782 84204
rect 258902 84192 258908 84204
rect 258960 84192 258966 84244
rect 244458 84164 244464 84176
rect 244419 84136 244464 84164
rect 244458 84124 244464 84136
rect 244516 84124 244522 84176
rect 245010 84124 245016 84176
rect 245068 84164 245074 84176
rect 245102 84164 245108 84176
rect 245068 84136 245108 84164
rect 245068 84124 245074 84136
rect 245102 84124 245108 84136
rect 245160 84124 245166 84176
rect 261662 84164 261668 84176
rect 261623 84136 261668 84164
rect 261662 84124 261668 84136
rect 261720 84124 261726 84176
rect 264514 84164 264520 84176
rect 264475 84136 264520 84164
rect 264514 84124 264520 84136
rect 264572 84124 264578 84176
rect 265802 84124 265808 84176
rect 265860 84164 265866 84176
rect 266354 84164 266360 84176
rect 265860 84136 266360 84164
rect 265860 84124 265866 84136
rect 266354 84124 266360 84136
rect 266412 84124 266418 84176
rect 293310 84164 293316 84176
rect 293271 84136 293316 84164
rect 293310 84124 293316 84136
rect 293368 84124 293374 84176
rect 294782 84164 294788 84176
rect 294743 84136 294788 84164
rect 294782 84124 294788 84136
rect 294840 84124 294846 84176
rect 319622 84164 319628 84176
rect 319583 84136 319628 84164
rect 319622 84124 319628 84136
rect 319680 84124 319686 84176
rect 326246 84124 326252 84176
rect 326304 84164 326310 84176
rect 326338 84164 326344 84176
rect 326304 84136 326344 84164
rect 326304 84124 326310 84136
rect 326338 84124 326344 84136
rect 326396 84124 326402 84176
rect 253014 84056 253020 84108
rect 253072 84096 253078 84108
rect 253106 84096 253112 84108
rect 253072 84068 253112 84096
rect 253072 84056 253078 84068
rect 253106 84056 253112 84068
rect 253164 84056 253170 84108
rect 263042 83008 263048 83020
rect 263003 82980 263048 83008
rect 263042 82968 263048 82980
rect 263100 82968 263106 83020
rect 320818 82940 320824 82952
rect 320779 82912 320824 82940
rect 320818 82900 320824 82912
rect 320876 82900 320882 82952
rect 320818 82804 320824 82816
rect 320779 82776 320824 82804
rect 320818 82764 320824 82776
rect 320876 82764 320882 82816
rect 329009 82807 329067 82813
rect 329009 82773 329021 82807
rect 329055 82804 329067 82807
rect 329190 82804 329196 82816
rect 329055 82776 329196 82804
rect 329055 82773 329067 82776
rect 329009 82767 329067 82773
rect 329190 82764 329196 82776
rect 329248 82764 329254 82816
rect 232038 81404 232044 81456
rect 232096 81444 232102 81456
rect 232130 81444 232136 81456
rect 232096 81416 232136 81444
rect 232096 81404 232102 81416
rect 232130 81404 232136 81416
rect 232188 81404 232194 81456
rect 231210 80112 231216 80164
rect 231268 80112 231274 80164
rect 243630 80152 243636 80164
rect 243556 80124 243636 80152
rect 231228 80028 231256 80112
rect 243556 80028 243584 80124
rect 243630 80112 243636 80124
rect 243688 80112 243694 80164
rect 231210 79976 231216 80028
rect 231268 79976 231274 80028
rect 243538 79976 243544 80028
rect 243596 79976 243602 80028
rect 246025 77367 246083 77373
rect 246025 77333 246037 77367
rect 246071 77364 246083 77367
rect 246114 77364 246120 77376
rect 246071 77336 246120 77364
rect 246071 77333 246083 77336
rect 246025 77327 246083 77333
rect 246114 77324 246120 77336
rect 246172 77324 246178 77376
rect 100662 77228 100668 77240
rect 100623 77200 100668 77228
rect 100662 77188 100668 77200
rect 100720 77188 100726 77240
rect 243538 77188 243544 77240
rect 243596 77228 243602 77240
rect 243630 77228 243636 77240
rect 243596 77200 243636 77228
rect 243596 77188 243602 77200
rect 243630 77188 243636 77200
rect 243688 77188 243694 77240
rect 244458 77228 244464 77240
rect 244419 77200 244464 77228
rect 244458 77188 244464 77200
rect 244516 77188 244522 77240
rect 314194 77228 314200 77240
rect 314155 77200 314200 77228
rect 314194 77188 314200 77200
rect 314252 77188 314258 77240
rect 317046 77188 317052 77240
rect 317104 77188 317110 77240
rect 318153 77231 318211 77237
rect 318153 77197 318165 77231
rect 318199 77228 318211 77231
rect 318242 77228 318248 77240
rect 318199 77200 318248 77228
rect 318199 77197 318211 77200
rect 318153 77191 318211 77197
rect 318242 77188 318248 77200
rect 318300 77188 318306 77240
rect 314378 77120 314384 77172
rect 314436 77120 314442 77172
rect 314396 77036 314424 77120
rect 317064 77104 317092 77188
rect 317046 77052 317052 77104
rect 317104 77052 317110 77104
rect 314378 76984 314384 77036
rect 314436 76984 314442 77036
rect 258902 76004 258908 76016
rect 258828 75976 258908 76004
rect 107470 75936 107476 75948
rect 107431 75908 107476 75936
rect 107470 75896 107476 75908
rect 107528 75896 107534 75948
rect 232317 75939 232375 75945
rect 232317 75905 232329 75939
rect 232363 75936 232375 75939
rect 232406 75936 232412 75948
rect 232363 75908 232412 75936
rect 232363 75905 232375 75908
rect 232317 75899 232375 75905
rect 232406 75896 232412 75908
rect 232464 75896 232470 75948
rect 258828 75880 258856 75976
rect 258902 75964 258908 75976
rect 258960 75964 258966 76016
rect 260374 76004 260380 76016
rect 260300 75976 260380 76004
rect 260300 75880 260328 75976
rect 260374 75964 260380 75976
rect 260432 75964 260438 76016
rect 333146 75964 333152 76016
rect 333204 75964 333210 76016
rect 331766 75896 331772 75948
rect 331824 75896 331830 75948
rect 254762 75868 254768 75880
rect 254723 75840 254768 75868
rect 254762 75828 254768 75840
rect 254820 75828 254826 75880
rect 258810 75828 258816 75880
rect 258868 75828 258874 75880
rect 260282 75828 260288 75880
rect 260340 75828 260346 75880
rect 331784 75868 331812 75896
rect 333164 75880 333192 75964
rect 333238 75896 333244 75948
rect 333296 75896 333302 75948
rect 341426 75896 341432 75948
rect 341484 75936 341490 75948
rect 341702 75936 341708 75948
rect 341484 75908 341708 75936
rect 341484 75896 341490 75908
rect 341702 75896 341708 75908
rect 341760 75896 341766 75948
rect 331858 75868 331864 75880
rect 331784 75840 331864 75868
rect 331858 75828 331864 75840
rect 331916 75828 331922 75880
rect 333146 75828 333152 75880
rect 333204 75828 333210 75880
rect 333256 75868 333284 75896
rect 333330 75868 333336 75880
rect 333256 75840 333336 75868
rect 333330 75828 333336 75840
rect 333388 75828 333394 75880
rect 322290 74740 322296 74792
rect 322348 74740 322354 74792
rect 322308 74656 322336 74740
rect 261662 74644 261668 74656
rect 261623 74616 261668 74644
rect 261662 74604 261668 74616
rect 261720 74604 261726 74656
rect 322290 74604 322296 74656
rect 322348 74604 322354 74656
rect 246022 74576 246028 74588
rect 245983 74548 246028 74576
rect 246022 74536 246028 74548
rect 246080 74536 246086 74588
rect 253106 74536 253112 74588
rect 253164 74536 253170 74588
rect 257062 74536 257068 74588
rect 257120 74576 257126 74588
rect 257154 74576 257160 74588
rect 257120 74548 257160 74576
rect 257120 74536 257126 74548
rect 257154 74536 257160 74548
rect 257212 74536 257218 74588
rect 264514 74536 264520 74588
rect 264572 74576 264578 74588
rect 293310 74576 293316 74588
rect 264572 74548 264617 74576
rect 293271 74548 293316 74576
rect 264572 74536 264578 74548
rect 293310 74536 293316 74548
rect 293368 74536 293374 74588
rect 294782 74576 294788 74588
rect 294743 74548 294788 74576
rect 294782 74536 294788 74548
rect 294840 74536 294846 74588
rect 295978 74536 295984 74588
rect 296036 74576 296042 74588
rect 296070 74576 296076 74588
rect 296036 74548 296076 74576
rect 296036 74536 296042 74548
rect 296070 74536 296076 74548
rect 296128 74536 296134 74588
rect 319622 74576 319628 74588
rect 319583 74548 319628 74576
rect 319622 74536 319628 74548
rect 319680 74536 319686 74588
rect 253124 74440 253152 74536
rect 265618 74468 265624 74520
rect 265676 74508 265682 74520
rect 265802 74508 265808 74520
rect 265676 74480 265808 74508
rect 265676 74468 265682 74480
rect 265802 74468 265808 74480
rect 265860 74468 265866 74520
rect 322290 74468 322296 74520
rect 322348 74468 322354 74520
rect 253290 74440 253296 74452
rect 253124 74412 253296 74440
rect 253290 74400 253296 74412
rect 253348 74400 253354 74452
rect 322308 74440 322336 74468
rect 322382 74440 322388 74452
rect 322308 74412 322388 74440
rect 322382 74400 322388 74412
rect 322440 74400 322446 74452
rect 320821 73219 320879 73225
rect 320821 73185 320833 73219
rect 320867 73216 320879 73219
rect 321094 73216 321100 73228
rect 320867 73188 321100 73216
rect 320867 73185 320879 73188
rect 320821 73179 320879 73185
rect 321094 73176 321100 73188
rect 321152 73176 321158 73228
rect 253201 73151 253259 73157
rect 253201 73117 253213 73151
rect 253247 73148 253259 73151
rect 253290 73148 253296 73160
rect 253247 73120 253296 73148
rect 253247 73117 253259 73120
rect 253201 73111 253259 73117
rect 253290 73108 253296 73120
rect 253348 73108 253354 73160
rect 232130 73080 232136 73092
rect 232091 73052 232136 73080
rect 232130 73040 232136 73052
rect 232188 73040 232194 73092
rect 329006 71788 329012 71800
rect 328967 71760 329012 71788
rect 329006 71748 329012 71760
rect 329064 71748 329070 71800
rect 254765 69683 254823 69689
rect 254765 69649 254777 69683
rect 254811 69680 254823 69683
rect 254946 69680 254952 69692
rect 254811 69652 254952 69680
rect 254811 69649 254823 69652
rect 254765 69643 254823 69649
rect 254946 69640 254952 69652
rect 255004 69640 255010 69692
rect 100662 67640 100668 67652
rect 100623 67612 100668 67640
rect 100662 67600 100668 67612
rect 100720 67600 100726 67652
rect 231118 67600 231124 67652
rect 231176 67640 231182 67652
rect 231302 67640 231308 67652
rect 231176 67612 231308 67640
rect 231176 67600 231182 67612
rect 231302 67600 231308 67612
rect 231360 67600 231366 67652
rect 232590 67600 232596 67652
rect 232648 67640 232654 67652
rect 232682 67640 232688 67652
rect 232648 67612 232688 67640
rect 232648 67600 232654 67612
rect 232682 67600 232688 67612
rect 232740 67600 232746 67652
rect 263042 67640 263048 67652
rect 263003 67612 263048 67640
rect 263042 67600 263048 67612
rect 263100 67600 263106 67652
rect 314194 67640 314200 67652
rect 314155 67612 314200 67640
rect 314194 67600 314200 67612
rect 314252 67600 314258 67652
rect 316862 67600 316868 67652
rect 316920 67640 316926 67652
rect 316954 67640 316960 67652
rect 316920 67612 316960 67640
rect 316920 67600 316926 67612
rect 316954 67600 316960 67612
rect 317012 67600 317018 67652
rect 318150 67640 318156 67652
rect 318111 67612 318156 67640
rect 318150 67600 318156 67612
rect 318208 67600 318214 67652
rect 345382 67572 345388 67584
rect 345343 67544 345388 67572
rect 345382 67532 345388 67544
rect 345440 67532 345446 67584
rect 260282 66348 260288 66360
rect 260208 66320 260288 66348
rect 260208 66292 260236 66320
rect 260282 66308 260288 66320
rect 260340 66308 260346 66360
rect 260190 66240 260196 66292
rect 260248 66240 260254 66292
rect 330386 66240 330392 66292
rect 330444 66280 330450 66292
rect 330478 66280 330484 66292
rect 330444 66252 330484 66280
rect 330444 66240 330450 66252
rect 330478 66240 330484 66252
rect 330536 66240 330542 66292
rect 331766 66240 331772 66292
rect 331824 66280 331830 66292
rect 331858 66280 331864 66292
rect 331824 66252 331864 66280
rect 331824 66240 331830 66252
rect 331858 66240 331864 66252
rect 331916 66240 331922 66292
rect 333238 66240 333244 66292
rect 333296 66280 333302 66292
rect 333330 66280 333336 66292
rect 333296 66252 333336 66280
rect 333296 66240 333302 66252
rect 333330 66240 333336 66252
rect 333388 66240 333394 66292
rect 334526 66240 334532 66292
rect 334584 66280 334590 66292
rect 334618 66280 334624 66292
rect 334584 66252 334624 66280
rect 334584 66240 334590 66252
rect 334618 66240 334624 66252
rect 334676 66240 334682 66292
rect 335814 66240 335820 66292
rect 335872 66280 335878 66292
rect 335906 66280 335912 66292
rect 335872 66252 335912 66280
rect 335872 66240 335878 66252
rect 335906 66240 335912 66252
rect 335964 66240 335970 66292
rect 107470 66212 107476 66224
rect 107431 66184 107476 66212
rect 107470 66172 107476 66184
rect 107528 66172 107534 66224
rect 231118 66172 231124 66224
rect 231176 66212 231182 66224
rect 231302 66212 231308 66224
rect 231176 66184 231308 66212
rect 231176 66172 231182 66184
rect 231302 66172 231308 66184
rect 231360 66172 231366 66224
rect 232314 66172 232320 66224
rect 232372 66212 232378 66224
rect 232406 66212 232412 66224
rect 232372 66184 232412 66212
rect 232372 66172 232378 66184
rect 232406 66172 232412 66184
rect 232464 66172 232470 66224
rect 314194 66212 314200 66224
rect 314155 66184 314200 66212
rect 314194 66172 314200 66184
rect 314252 66172 314258 66224
rect 258810 64880 258816 64932
rect 258868 64920 258874 64932
rect 258902 64920 258908 64932
rect 258868 64892 258908 64920
rect 258868 64880 258874 64892
rect 258902 64880 258908 64892
rect 258960 64880 258966 64932
rect 260190 64812 260196 64864
rect 260248 64852 260254 64864
rect 260374 64852 260380 64864
rect 260248 64824 260380 64852
rect 260248 64812 260254 64824
rect 260374 64812 260380 64824
rect 260432 64812 260438 64864
rect 264514 64852 264520 64864
rect 264475 64824 264520 64852
rect 264514 64812 264520 64824
rect 264572 64812 264578 64864
rect 265802 64852 265808 64864
rect 265763 64824 265808 64852
rect 265802 64812 265808 64824
rect 265860 64812 265866 64864
rect 293310 64852 293316 64864
rect 293271 64824 293316 64852
rect 293310 64812 293316 64824
rect 293368 64812 293374 64864
rect 294782 64852 294788 64864
rect 294743 64824 294788 64852
rect 294782 64812 294788 64824
rect 294840 64812 294846 64864
rect 319622 64852 319628 64864
rect 319583 64824 319628 64852
rect 319622 64812 319628 64824
rect 319680 64812 319686 64864
rect 322293 64855 322351 64861
rect 322293 64821 322305 64855
rect 322339 64852 322351 64855
rect 322382 64852 322388 64864
rect 322339 64824 322388 64852
rect 322339 64821 322351 64824
rect 322293 64815 322351 64821
rect 322382 64812 322388 64824
rect 322440 64812 322446 64864
rect 253198 63560 253204 63572
rect 253159 63532 253204 63560
rect 253198 63520 253204 63532
rect 253256 63520 253262 63572
rect 254765 63495 254823 63501
rect 254765 63461 254777 63495
rect 254811 63492 254823 63495
rect 254854 63492 254860 63504
rect 254811 63464 254860 63492
rect 254811 63461 254823 63464
rect 254765 63455 254823 63461
rect 254854 63452 254860 63464
rect 254912 63452 254918 63504
rect 321002 63492 321008 63504
rect 320963 63464 321008 63492
rect 321002 63452 321008 63464
rect 321060 63452 321066 63504
rect 326246 63452 326252 63504
rect 326304 63492 326310 63504
rect 326338 63492 326344 63504
rect 326304 63464 326344 63492
rect 326304 63452 326310 63464
rect 326338 63452 326344 63464
rect 326396 63452 326402 63504
rect 331766 63492 331772 63504
rect 331727 63464 331772 63492
rect 331766 63452 331772 63464
rect 331824 63452 331830 63504
rect 334526 61452 334532 61464
rect 334487 61424 334532 61452
rect 334526 61412 334532 61424
rect 334584 61412 334590 61464
rect 258902 60120 258908 60172
rect 258960 60120 258966 60172
rect 258920 60036 258948 60120
rect 258902 59984 258908 60036
rect 258960 59984 258966 60036
rect 296073 60027 296131 60033
rect 296073 59993 296085 60027
rect 296119 60024 296131 60027
rect 296162 60024 296168 60036
rect 296119 59996 296168 60024
rect 296119 59993 296131 59996
rect 296073 59987 296131 59993
rect 296162 59984 296168 59996
rect 296220 59984 296226 60036
rect 244918 57944 244924 57996
rect 244976 57984 244982 57996
rect 245010 57984 245016 57996
rect 244976 57956 245016 57984
rect 244976 57944 244982 57956
rect 245010 57944 245016 57956
rect 245068 57944 245074 57996
rect 345382 57984 345388 57996
rect 345343 57956 345388 57984
rect 345382 57944 345388 57956
rect 345440 57944 345446 57996
rect 100662 57916 100668 57928
rect 100623 57888 100668 57916
rect 100662 57876 100668 57888
rect 100720 57876 100726 57928
rect 246485 57919 246543 57925
rect 246485 57885 246497 57919
rect 246531 57916 246543 57919
rect 246574 57916 246580 57928
rect 246531 57888 246580 57916
rect 246531 57885 246543 57888
rect 246485 57879 246543 57885
rect 246574 57876 246580 57888
rect 246632 57876 246638 57928
rect 107470 56624 107476 56636
rect 107431 56596 107476 56624
rect 107470 56584 107476 56596
rect 107528 56584 107534 56636
rect 314194 56624 314200 56636
rect 314155 56596 314200 56624
rect 314194 56584 314200 56596
rect 314252 56584 314258 56636
rect 240597 56559 240655 56565
rect 240597 56525 240609 56559
rect 240643 56556 240655 56559
rect 240686 56556 240692 56568
rect 240643 56528 240692 56556
rect 240643 56525 240655 56528
rect 240597 56519 240655 56525
rect 240686 56516 240692 56528
rect 240744 56516 240750 56568
rect 244458 56516 244464 56568
rect 244516 56556 244522 56568
rect 244516 56528 244561 56556
rect 244516 56516 244522 56528
rect 261573 56015 261631 56021
rect 261573 55981 261585 56015
rect 261619 56012 261631 56015
rect 261662 56012 261668 56024
rect 261619 55984 261668 56012
rect 261619 55981 261631 55984
rect 261573 55975 261631 55981
rect 261662 55972 261668 55984
rect 261720 55972 261726 56024
rect 265802 55332 265808 55344
rect 265763 55304 265808 55332
rect 265802 55292 265808 55304
rect 265860 55292 265866 55344
rect 322290 55332 322296 55344
rect 322251 55304 322296 55332
rect 322290 55292 322296 55304
rect 322348 55292 322354 55344
rect 231302 55196 231308 55208
rect 231263 55168 231308 55196
rect 231302 55156 231308 55168
rect 231360 55156 231366 55208
rect 265802 55196 265808 55208
rect 265763 55168 265808 55196
rect 265802 55156 265808 55168
rect 265860 55156 265866 55208
rect 299014 55196 299020 55208
rect 298975 55168 299020 55196
rect 299014 55156 299020 55168
rect 299072 55156 299078 55208
rect 300302 55196 300308 55208
rect 300263 55168 300308 55196
rect 300302 55156 300308 55168
rect 300360 55156 300366 55208
rect 301774 55196 301780 55208
rect 301735 55168 301780 55196
rect 301774 55156 301780 55168
rect 301832 55156 301838 55208
rect 322290 55156 322296 55208
rect 322348 55196 322354 55208
rect 322382 55196 322388 55208
rect 322348 55168 322388 55196
rect 322348 55156 322354 55168
rect 322382 55156 322388 55168
rect 322440 55156 322446 55208
rect 254762 53836 254768 53848
rect 254723 53808 254768 53836
rect 254762 53796 254768 53808
rect 254820 53796 254826 53848
rect 331766 53836 331772 53848
rect 331727 53808 331772 53836
rect 331766 53796 331772 53808
rect 331824 53796 331830 53848
rect 326154 52436 326160 52488
rect 326212 52476 326218 52488
rect 326246 52476 326252 52488
rect 326212 52448 326252 52476
rect 326212 52436 326218 52448
rect 326246 52436 326252 52448
rect 326304 52436 326310 52488
rect 329006 52436 329012 52488
rect 329064 52476 329070 52488
rect 329190 52476 329196 52488
rect 329064 52448 329196 52476
rect 329064 52436 329070 52448
rect 329190 52436 329196 52448
rect 329248 52436 329254 52488
rect 333054 51076 333060 51128
rect 333112 51076 333118 51128
rect 333072 50980 333100 51076
rect 340046 51008 340052 51060
rect 340104 51048 340110 51060
rect 340230 51048 340236 51060
rect 340104 51020 340236 51048
rect 340104 51008 340110 51020
rect 340230 51008 340236 51020
rect 340288 51008 340294 51060
rect 333146 50980 333152 50992
rect 333072 50952 333152 50980
rect 333146 50940 333152 50952
rect 333204 50940 333210 50992
rect 253014 50328 253020 50380
rect 253072 50368 253078 50380
rect 253290 50368 253296 50380
rect 253072 50340 253296 50368
rect 253072 50328 253078 50340
rect 253290 50328 253296 50340
rect 253348 50328 253354 50380
rect 345382 48396 345388 48408
rect 345308 48368 345388 48396
rect 345308 48340 345336 48368
rect 345382 48356 345388 48368
rect 345440 48356 345446 48408
rect 100662 48328 100668 48340
rect 100623 48300 100668 48328
rect 100662 48288 100668 48300
rect 100720 48288 100726 48340
rect 244918 48288 244924 48340
rect 244976 48328 244982 48340
rect 245010 48328 245016 48340
rect 244976 48300 245016 48328
rect 244976 48288 244982 48300
rect 245010 48288 245016 48300
rect 245068 48288 245074 48340
rect 246482 48328 246488 48340
rect 246443 48300 246488 48328
rect 246482 48288 246488 48300
rect 246540 48288 246546 48340
rect 344186 48288 344192 48340
rect 344244 48328 344250 48340
rect 344278 48328 344284 48340
rect 344244 48300 344284 48328
rect 344244 48288 344250 48300
rect 344278 48288 344284 48300
rect 344336 48288 344342 48340
rect 345290 48288 345296 48340
rect 345348 48288 345354 48340
rect 257154 47064 257160 47116
rect 257212 47064 257218 47116
rect 240597 47039 240655 47045
rect 240597 47005 240609 47039
rect 240643 47036 240655 47039
rect 240686 47036 240692 47048
rect 240643 47008 240692 47036
rect 240643 47005 240655 47008
rect 240597 46999 240655 47005
rect 240686 46996 240692 47008
rect 240744 46996 240750 47048
rect 257172 46980 257200 47064
rect 232130 46968 232136 46980
rect 232091 46940 232136 46968
rect 232130 46928 232136 46940
rect 232188 46928 232194 46980
rect 244366 46928 244372 46980
rect 244424 46968 244430 46980
rect 244461 46971 244519 46977
rect 244461 46968 244473 46971
rect 244424 46940 244473 46968
rect 244424 46928 244430 46940
rect 244461 46937 244473 46940
rect 244507 46937 244519 46971
rect 244461 46931 244519 46937
rect 257154 46928 257160 46980
rect 257212 46928 257218 46980
rect 261570 46968 261576 46980
rect 261531 46940 261576 46968
rect 261570 46928 261576 46940
rect 261628 46928 261634 46980
rect 264514 46968 264520 46980
rect 264475 46940 264520 46968
rect 264514 46928 264520 46940
rect 264572 46928 264578 46980
rect 293313 46971 293371 46977
rect 293313 46937 293325 46971
rect 293359 46968 293371 46971
rect 293402 46968 293408 46980
rect 293359 46940 293408 46968
rect 293359 46937 293371 46940
rect 293313 46931 293371 46937
rect 293402 46928 293408 46940
rect 293460 46928 293466 46980
rect 294785 46971 294843 46977
rect 294785 46937 294797 46971
rect 294831 46968 294843 46971
rect 294874 46968 294880 46980
rect 294831 46940 294880 46968
rect 294831 46937 294843 46940
rect 294785 46931 294843 46937
rect 294874 46928 294880 46940
rect 294932 46928 294938 46980
rect 296073 46971 296131 46977
rect 296073 46937 296085 46971
rect 296119 46968 296131 46971
rect 296162 46968 296168 46980
rect 296119 46940 296168 46968
rect 296119 46937 296131 46940
rect 296073 46931 296131 46937
rect 296162 46928 296168 46940
rect 296220 46928 296226 46980
rect 319622 46968 319628 46980
rect 319583 46940 319628 46968
rect 319622 46928 319628 46940
rect 319680 46928 319686 46980
rect 334526 46968 334532 46980
rect 334487 46940 334532 46968
rect 334526 46928 334532 46940
rect 334584 46928 334590 46980
rect 341518 46928 341524 46980
rect 341576 46968 341582 46980
rect 341702 46968 341708 46980
rect 341576 46940 341708 46968
rect 341576 46928 341582 46940
rect 341702 46928 341708 46940
rect 341760 46928 341766 46980
rect 107470 46900 107476 46912
rect 107431 46872 107476 46900
rect 107470 46860 107476 46872
rect 107528 46860 107534 46912
rect 240686 46900 240692 46912
rect 240647 46872 240692 46900
rect 240686 46860 240692 46872
rect 240744 46860 240750 46912
rect 314194 46900 314200 46912
rect 314155 46872 314200 46900
rect 314194 46860 314200 46872
rect 314252 46860 314258 46912
rect 231302 45608 231308 45620
rect 231263 45580 231308 45608
rect 231302 45568 231308 45580
rect 231360 45568 231366 45620
rect 265802 45608 265808 45620
rect 265763 45580 265808 45608
rect 265802 45568 265808 45580
rect 265860 45568 265866 45620
rect 299014 45608 299020 45620
rect 298975 45580 299020 45608
rect 299014 45568 299020 45580
rect 299072 45568 299078 45620
rect 300302 45608 300308 45620
rect 300263 45580 300308 45608
rect 300302 45568 300308 45580
rect 300360 45568 300366 45620
rect 301774 45608 301780 45620
rect 301735 45580 301780 45608
rect 301774 45568 301780 45580
rect 301832 45568 301838 45620
rect 321005 45611 321063 45617
rect 321005 45577 321017 45611
rect 321051 45608 321063 45611
rect 321094 45608 321100 45620
rect 321051 45580 321100 45608
rect 321051 45577 321063 45580
rect 321005 45571 321063 45577
rect 321094 45568 321100 45580
rect 321152 45568 321158 45620
rect 252925 45543 252983 45549
rect 252925 45509 252937 45543
rect 252971 45540 252983 45543
rect 253014 45540 253020 45552
rect 252971 45512 253020 45540
rect 252971 45509 252983 45512
rect 252925 45503 252983 45509
rect 253014 45500 253020 45512
rect 253072 45500 253078 45552
rect 254762 45500 254768 45552
rect 254820 45500 254826 45552
rect 257154 45540 257160 45552
rect 257115 45512 257160 45540
rect 257154 45500 257160 45512
rect 257212 45500 257218 45552
rect 264425 45543 264483 45549
rect 264425 45509 264437 45543
rect 264471 45540 264483 45543
rect 264514 45540 264520 45552
rect 264471 45512 264520 45540
rect 264471 45509 264483 45512
rect 264425 45503 264483 45509
rect 264514 45500 264520 45512
rect 264572 45500 264578 45552
rect 319622 45540 319628 45552
rect 319583 45512 319628 45540
rect 319622 45500 319628 45512
rect 319680 45500 319686 45552
rect 322293 45543 322351 45549
rect 322293 45509 322305 45543
rect 322339 45540 322351 45543
rect 322382 45540 322388 45552
rect 322339 45512 322388 45540
rect 322339 45509 322351 45512
rect 322293 45503 322351 45509
rect 322382 45500 322388 45512
rect 322440 45500 322446 45552
rect 254780 45416 254808 45500
rect 254762 45364 254768 45416
rect 254820 45364 254826 45416
rect 326154 44208 326160 44260
rect 326212 44248 326218 44260
rect 326246 44248 326252 44260
rect 326212 44220 326252 44248
rect 326212 44208 326218 44220
rect 326246 44208 326252 44220
rect 326304 44208 326310 44260
rect 329006 44140 329012 44192
rect 329064 44180 329070 44192
rect 329098 44180 329104 44192
rect 329064 44152 329104 44180
rect 329064 44140 329070 44152
rect 329098 44140 329104 44152
rect 329156 44140 329162 44192
rect 326246 44072 326252 44124
rect 326304 44112 326310 44124
rect 326341 44115 326399 44121
rect 326341 44112 326353 44115
rect 326304 44084 326353 44112
rect 326304 44072 326310 44084
rect 326341 44081 326353 44084
rect 326387 44081 326399 44115
rect 326341 44075 326399 44081
rect 331766 44072 331772 44124
rect 331824 44112 331830 44124
rect 331950 44112 331956 44124
rect 331824 44084 331956 44112
rect 331824 44072 331830 44084
rect 331950 44072 331956 44084
rect 332008 44072 332014 44124
rect 261570 42140 261576 42152
rect 261531 42112 261576 42140
rect 261570 42100 261576 42112
rect 261628 42100 261634 42152
rect 244366 41460 244372 41472
rect 244327 41432 244372 41460
rect 244366 41420 244372 41432
rect 244424 41420 244430 41472
rect 344186 41460 344192 41472
rect 344112 41432 344192 41460
rect 344112 41404 344140 41432
rect 344186 41420 344192 41432
rect 344244 41420 344250 41472
rect 344094 41352 344100 41404
rect 344152 41352 344158 41404
rect 232317 40715 232375 40721
rect 232317 40681 232329 40715
rect 232363 40712 232375 40715
rect 232406 40712 232412 40724
rect 232363 40684 232412 40712
rect 232363 40681 232375 40684
rect 232317 40675 232375 40681
rect 232406 40672 232412 40684
rect 232464 40672 232470 40724
rect 232774 40712 232780 40724
rect 232735 40684 232780 40712
rect 232774 40672 232780 40684
rect 232832 40672 232838 40724
rect 252922 40712 252928 40724
rect 252883 40684 252928 40712
rect 252922 40672 252928 40684
rect 252980 40672 252986 40724
rect 321002 40712 321008 40724
rect 320963 40684 321008 40712
rect 321002 40672 321008 40684
rect 321060 40672 321066 40724
rect 322290 40712 322296 40724
rect 322251 40684 322296 40712
rect 322290 40672 322296 40684
rect 322348 40672 322354 40724
rect 335446 40264 335452 40316
rect 335504 40304 335510 40316
rect 344922 40304 344928 40316
rect 335504 40276 344928 40304
rect 335504 40264 335510 40276
rect 344922 40264 344928 40276
rect 344980 40264 344986 40316
rect 345290 38632 345296 38684
rect 345348 38672 345354 38684
rect 345382 38672 345388 38684
rect 345348 38644 345388 38672
rect 345348 38632 345354 38644
rect 345382 38632 345388 38644
rect 345440 38632 345446 38684
rect 100662 38604 100668 38616
rect 100623 38576 100668 38604
rect 100662 38564 100668 38576
rect 100720 38564 100726 38616
rect 244366 38604 244372 38616
rect 244327 38576 244372 38604
rect 244366 38564 244372 38576
rect 244424 38564 244430 38616
rect 240686 37380 240692 37392
rect 240647 37352 240692 37380
rect 240686 37340 240692 37352
rect 240744 37340 240750 37392
rect 265713 37383 265771 37389
rect 265713 37349 265725 37383
rect 265759 37380 265771 37383
rect 265802 37380 265808 37392
rect 265759 37352 265808 37380
rect 265759 37349 265771 37352
rect 265713 37343 265771 37349
rect 265802 37340 265808 37352
rect 265860 37340 265866 37392
rect 107470 37312 107476 37324
rect 107431 37284 107476 37312
rect 107470 37272 107476 37284
rect 107528 37272 107534 37324
rect 258810 37272 258816 37324
rect 258868 37312 258874 37324
rect 258902 37312 258908 37324
rect 258868 37284 258908 37312
rect 258868 37272 258874 37284
rect 258902 37272 258908 37284
rect 258960 37272 258966 37324
rect 314194 37312 314200 37324
rect 314155 37284 314200 37312
rect 314194 37272 314200 37284
rect 314252 37272 314258 37324
rect 240226 37204 240232 37256
rect 240284 37244 240290 37256
rect 240686 37244 240692 37256
rect 240284 37216 240692 37244
rect 240284 37204 240290 37216
rect 240686 37204 240692 37216
rect 240744 37204 240750 37256
rect 261573 35955 261631 35961
rect 261573 35921 261585 35955
rect 261619 35952 261631 35955
rect 261662 35952 261668 35964
rect 261619 35924 261668 35952
rect 261619 35921 261631 35924
rect 261573 35915 261631 35921
rect 261662 35912 261668 35924
rect 261720 35912 261726 35964
rect 264422 35952 264428 35964
rect 264383 35924 264428 35952
rect 264422 35912 264428 35924
rect 264480 35912 264486 35964
rect 265710 35952 265716 35964
rect 265671 35924 265716 35952
rect 265710 35912 265716 35924
rect 265768 35912 265774 35964
rect 319622 35952 319628 35964
rect 319583 35924 319628 35952
rect 319622 35912 319628 35924
rect 319680 35912 319686 35964
rect 252922 35884 252928 35896
rect 252883 35856 252928 35884
rect 252922 35844 252928 35856
rect 252980 35844 252986 35896
rect 299014 35884 299020 35896
rect 298975 35856 299020 35884
rect 299014 35844 299020 35856
rect 299072 35844 299078 35896
rect 300302 35884 300308 35896
rect 300263 35856 300308 35884
rect 300302 35844 300308 35856
rect 300360 35844 300366 35896
rect 301774 35884 301780 35896
rect 301735 35856 301780 35884
rect 301774 35844 301780 35856
rect 301832 35844 301838 35896
rect 245838 33804 245844 33856
rect 245896 33844 245902 33856
rect 246022 33844 246028 33856
rect 245896 33816 246028 33844
rect 245896 33804 245902 33816
rect 246022 33804 246028 33816
rect 246080 33804 246086 33856
rect 262950 31764 262956 31816
rect 263008 31764 263014 31816
rect 319622 31804 319628 31816
rect 319548 31776 319628 31804
rect 262968 31668 262996 31764
rect 319548 31748 319576 31776
rect 319622 31764 319628 31776
rect 319680 31764 319686 31816
rect 319530 31696 319536 31748
rect 319588 31696 319594 31748
rect 321002 31736 321008 31748
rect 320963 31708 321008 31736
rect 321002 31696 321008 31708
rect 321060 31696 321066 31748
rect 263042 31668 263048 31680
rect 262968 31640 263048 31668
rect 263042 31628 263048 31640
rect 263100 31628 263106 31680
rect 379422 29180 379428 29232
rect 379480 29220 379486 29232
rect 386322 29220 386328 29232
rect 379480 29192 386328 29220
rect 379480 29180 379486 29192
rect 386322 29180 386328 29192
rect 386380 29180 386386 29232
rect 240594 29044 240600 29096
rect 240652 29044 240658 29096
rect 100662 29016 100668 29028
rect 100623 28988 100668 29016
rect 100662 28976 100668 28988
rect 100720 28976 100726 29028
rect 240612 28960 240640 29044
rect 264422 28976 264428 29028
rect 264480 29016 264486 29028
rect 264514 29016 264520 29028
rect 264480 28988 264520 29016
rect 264480 28976 264486 28988
rect 264514 28976 264520 28988
rect 264572 28976 264578 29028
rect 265710 28976 265716 29028
rect 265768 29016 265774 29028
rect 265802 29016 265808 29028
rect 265768 28988 265808 29016
rect 265768 28976 265774 28988
rect 265802 28976 265808 28988
rect 265860 28976 265866 29028
rect 267090 28976 267096 29028
rect 267148 29016 267154 29028
rect 267182 29016 267188 29028
rect 267148 28988 267188 29016
rect 267148 28976 267154 28988
rect 267182 28976 267188 28988
rect 267240 28976 267246 29028
rect 268562 28976 268568 29028
rect 268620 29016 268626 29028
rect 268654 29016 268660 29028
rect 268620 28988 268660 29016
rect 268620 28976 268626 28988
rect 268654 28976 268660 28988
rect 268712 28976 268718 29028
rect 333054 28976 333060 29028
rect 333112 28976 333118 29028
rect 240594 28908 240600 28960
rect 240652 28908 240658 28960
rect 244918 28908 244924 28960
rect 244976 28948 244982 28960
rect 245010 28948 245016 28960
rect 244976 28920 245016 28948
rect 244976 28908 244982 28920
rect 245010 28908 245016 28920
rect 245068 28908 245074 28960
rect 333072 28880 333100 28976
rect 340046 28948 340052 28960
rect 339972 28920 340052 28948
rect 339972 28892 340000 28920
rect 340046 28908 340052 28920
rect 340104 28908 340110 28960
rect 333146 28880 333152 28892
rect 333072 28852 333152 28880
rect 333146 28840 333152 28852
rect 333204 28840 333210 28892
rect 339954 28840 339960 28892
rect 340012 28840 340018 28892
rect 232314 27656 232320 27668
rect 232275 27628 232320 27656
rect 232314 27616 232320 27628
rect 232372 27616 232378 27668
rect 232774 27656 232780 27668
rect 232735 27628 232780 27656
rect 232774 27616 232780 27628
rect 232832 27616 232838 27668
rect 257154 27656 257160 27668
rect 257115 27628 257160 27656
rect 257154 27616 257160 27628
rect 257212 27616 257218 27668
rect 326338 27656 326344 27668
rect 326299 27628 326344 27656
rect 326338 27616 326344 27628
rect 326396 27616 326402 27668
rect 107470 27588 107476 27600
rect 107431 27560 107476 27588
rect 107470 27548 107476 27560
rect 107528 27548 107534 27600
rect 244458 27588 244464 27600
rect 244419 27560 244464 27588
rect 244458 27548 244464 27560
rect 244516 27548 244522 27600
rect 314194 27588 314200 27600
rect 314155 27560 314200 27588
rect 314194 27548 314200 27560
rect 314252 27548 314258 27600
rect 252925 26299 252983 26305
rect 252925 26265 252937 26299
rect 252971 26296 252983 26299
rect 253014 26296 253020 26308
rect 252971 26268 253020 26296
rect 252971 26265 252983 26268
rect 252925 26259 252983 26265
rect 253014 26256 253020 26268
rect 253072 26256 253078 26308
rect 299014 26296 299020 26308
rect 298975 26268 299020 26296
rect 299014 26256 299020 26268
rect 299072 26256 299078 26308
rect 300302 26296 300308 26308
rect 300263 26268 300308 26296
rect 300302 26256 300308 26268
rect 300360 26256 300366 26308
rect 301774 26296 301780 26308
rect 301735 26268 301780 26296
rect 301774 26256 301780 26268
rect 301832 26256 301838 26308
rect 329190 24828 329196 24880
rect 329248 24868 329254 24880
rect 329374 24868 329380 24880
rect 329248 24840 329380 24868
rect 329248 24828 329254 24840
rect 329374 24828 329380 24840
rect 329432 24828 329438 24880
rect 297634 23400 297640 23452
rect 297692 23440 297698 23452
rect 300673 23443 300731 23449
rect 300673 23440 300685 23443
rect 297692 23412 300685 23440
rect 297692 23400 297698 23412
rect 300673 23409 300685 23412
rect 300719 23409 300731 23443
rect 300673 23403 300731 23409
rect 297542 23372 297548 23384
rect 297503 23344 297548 23372
rect 297542 23332 297548 23344
rect 297600 23332 297606 23384
rect 2866 22040 2872 22092
rect 2924 22080 2930 22092
rect 349798 22080 349804 22092
rect 2924 22052 349804 22080
rect 2924 22040 2930 22052
rect 349798 22040 349804 22052
rect 349856 22040 349862 22092
rect 326338 19428 326344 19440
rect 326172 19400 326344 19428
rect 326172 19372 326200 19400
rect 326338 19388 326344 19400
rect 326396 19388 326402 19440
rect 237926 19320 237932 19372
rect 237984 19360 237990 19372
rect 238018 19360 238024 19372
rect 237984 19332 238024 19360
rect 237984 19320 237990 19332
rect 238018 19320 238024 19332
rect 238076 19320 238082 19372
rect 242158 19320 242164 19372
rect 242216 19360 242222 19372
rect 242250 19360 242256 19372
rect 242216 19332 242256 19360
rect 242216 19320 242222 19332
rect 242250 19320 242256 19332
rect 242308 19320 242314 19372
rect 243538 19320 243544 19372
rect 243596 19360 243602 19372
rect 243630 19360 243636 19372
rect 243596 19332 243636 19360
rect 243596 19320 243602 19332
rect 243630 19320 243636 19332
rect 243688 19320 243694 19372
rect 245838 19320 245844 19372
rect 245896 19360 245902 19372
rect 246022 19360 246028 19372
rect 245896 19332 246028 19360
rect 245896 19320 245902 19332
rect 246022 19320 246028 19332
rect 246080 19320 246086 19372
rect 326154 19320 326160 19372
rect 326212 19320 326218 19372
rect 344094 19320 344100 19372
rect 344152 19360 344158 19372
rect 344186 19360 344192 19372
rect 344152 19332 344192 19360
rect 344152 19320 344158 19332
rect 344186 19320 344192 19332
rect 344244 19320 344250 19372
rect 345382 19320 345388 19372
rect 345440 19360 345446 19372
rect 345474 19360 345480 19372
rect 345440 19332 345480 19360
rect 345440 19320 345446 19332
rect 345474 19320 345480 19332
rect 345532 19320 345538 19372
rect 100478 19252 100484 19304
rect 100536 19292 100542 19304
rect 100662 19292 100668 19304
rect 100536 19264 100668 19292
rect 100536 19252 100542 19264
rect 100662 19252 100668 19264
rect 100720 19252 100726 19304
rect 110322 19252 110328 19304
rect 110380 19292 110386 19304
rect 346578 19292 346584 19304
rect 110380 19264 346584 19292
rect 110380 19252 110386 19264
rect 346578 19252 346584 19264
rect 346636 19252 346642 19304
rect 103422 19184 103428 19236
rect 103480 19224 103486 19236
rect 345658 19224 345664 19236
rect 103480 19196 345664 19224
rect 103480 19184 103486 19196
rect 345658 19184 345664 19196
rect 345716 19184 345722 19236
rect 99282 19116 99288 19168
rect 99340 19156 99346 19168
rect 343910 19156 343916 19168
rect 99340 19128 343916 19156
rect 99340 19116 99346 19128
rect 343910 19116 343916 19128
rect 343968 19116 343974 19168
rect 96522 19048 96528 19100
rect 96580 19088 96586 19100
rect 342530 19088 342536 19100
rect 96580 19060 342536 19088
rect 96580 19048 96586 19060
rect 342530 19048 342536 19060
rect 342588 19048 342594 19100
rect 92382 18980 92388 19032
rect 92440 19020 92446 19032
rect 342806 19020 342812 19032
rect 92440 18992 342812 19020
rect 92440 18980 92446 18992
rect 342806 18980 342812 18992
rect 342864 18980 342870 19032
rect 89622 18912 89628 18964
rect 89680 18952 89686 18964
rect 341334 18952 341340 18964
rect 89680 18924 341340 18952
rect 89680 18912 89686 18924
rect 341334 18912 341340 18924
rect 341392 18912 341398 18964
rect 85482 18844 85488 18896
rect 85540 18884 85546 18896
rect 341058 18884 341064 18896
rect 85540 18856 341064 18884
rect 85540 18844 85546 18856
rect 341058 18844 341064 18856
rect 341116 18844 341122 18896
rect 82630 18776 82636 18828
rect 82688 18816 82694 18828
rect 339770 18816 339776 18828
rect 82688 18788 339776 18816
rect 82688 18776 82694 18788
rect 339770 18776 339776 18788
rect 339828 18776 339834 18828
rect 78582 18708 78588 18760
rect 78640 18748 78646 18760
rect 339862 18748 339868 18760
rect 78640 18720 339868 18748
rect 78640 18708 78646 18720
rect 339862 18708 339868 18720
rect 339920 18708 339926 18760
rect 74442 18640 74448 18692
rect 74500 18680 74506 18692
rect 338482 18680 338488 18692
rect 74500 18652 338488 18680
rect 74500 18640 74506 18652
rect 338482 18640 338488 18652
rect 338540 18640 338546 18692
rect 5442 18572 5448 18624
rect 5500 18612 5506 18624
rect 324866 18612 324872 18624
rect 5500 18584 324872 18612
rect 5500 18572 5506 18584
rect 324866 18572 324872 18584
rect 324924 18572 324930 18624
rect 294874 18504 294880 18556
rect 294932 18544 294938 18556
rect 442994 18544 443000 18556
rect 294932 18516 443000 18544
rect 294932 18504 294938 18516
rect 442994 18504 443000 18516
rect 443052 18504 443058 18556
rect 301774 18272 301780 18284
rect 301735 18244 301780 18272
rect 301774 18232 301780 18244
rect 301832 18232 301838 18284
rect 301866 18204 301872 18216
rect 301827 18176 301872 18204
rect 301866 18164 301872 18176
rect 301924 18164 301930 18216
rect 304629 18071 304687 18077
rect 304629 18037 304641 18071
rect 304675 18068 304687 18071
rect 304810 18068 304816 18080
rect 304675 18040 304816 18068
rect 304675 18037 304687 18040
rect 304629 18031 304687 18037
rect 304810 18028 304816 18040
rect 304868 18028 304874 18080
rect 322934 18028 322940 18080
rect 322992 18068 322998 18080
rect 332502 18068 332508 18080
rect 322992 18040 332508 18068
rect 322992 18028 322998 18040
rect 332502 18028 332508 18040
rect 332560 18028 332566 18080
rect 240226 17960 240232 18012
rect 240284 18000 240290 18012
rect 240686 18000 240692 18012
rect 240284 17972 240692 18000
rect 240284 17960 240290 17972
rect 240686 17960 240692 17972
rect 240744 17960 240750 18012
rect 244458 18000 244464 18012
rect 244419 17972 244464 18000
rect 244458 17960 244464 17972
rect 244516 17960 244522 18012
rect 246298 17960 246304 18012
rect 246356 18000 246362 18012
rect 246482 18000 246488 18012
rect 246356 17972 246488 18000
rect 246356 17960 246362 17972
rect 246482 17960 246488 17972
rect 246540 17960 246546 18012
rect 304902 18000 304908 18012
rect 304863 17972 304908 18000
rect 304902 17960 304908 17972
rect 304960 17960 304966 18012
rect 314194 18000 314200 18012
rect 314155 17972 314200 18000
rect 314194 17960 314200 17972
rect 314252 17960 314258 18012
rect 329098 18000 329104 18012
rect 329059 17972 329104 18000
rect 329098 17960 329104 17972
rect 329156 17960 329162 18012
rect 293678 17892 293684 17944
rect 293736 17932 293742 17944
rect 431954 17932 431960 17944
rect 293736 17904 431960 17932
rect 293736 17892 293742 17904
rect 431954 17892 431960 17904
rect 432012 17892 432018 17944
rect 253106 17824 253112 17876
rect 253164 17864 253170 17876
rect 253290 17864 253296 17876
rect 253164 17836 253296 17864
rect 253164 17824 253170 17836
rect 253290 17824 253296 17836
rect 253348 17824 253354 17876
rect 293402 17824 293408 17876
rect 293460 17864 293466 17876
rect 433334 17864 433340 17876
rect 293460 17836 433340 17864
rect 293460 17824 293466 17836
rect 433334 17824 433340 17836
rect 433392 17824 433398 17876
rect 293586 17756 293592 17808
rect 293644 17796 293650 17808
rect 434714 17796 434720 17808
rect 293644 17768 434720 17796
rect 293644 17756 293650 17768
rect 434714 17756 434720 17768
rect 434772 17756 434778 17808
rect 293494 17688 293500 17740
rect 293552 17728 293558 17740
rect 436094 17728 436100 17740
rect 293552 17700 436100 17728
rect 293552 17688 293558 17700
rect 436094 17688 436100 17700
rect 436152 17688 436158 17740
rect 294966 17620 294972 17672
rect 295024 17660 295030 17672
rect 438854 17660 438860 17672
rect 295024 17632 438860 17660
rect 295024 17620 295030 17632
rect 438854 17620 438860 17632
rect 438912 17620 438918 17672
rect 295058 17552 295064 17604
rect 295116 17592 295122 17604
rect 440234 17592 440240 17604
rect 295116 17564 440240 17592
rect 295116 17552 295122 17564
rect 440234 17552 440240 17564
rect 440292 17552 440298 17604
rect 303062 17484 303068 17536
rect 303120 17524 303126 17536
rect 483014 17524 483020 17536
rect 303120 17496 483020 17524
rect 303120 17484 303126 17496
rect 483014 17484 483020 17496
rect 483072 17484 483078 17536
rect 304626 17416 304632 17468
rect 304684 17456 304690 17468
rect 485774 17456 485780 17468
rect 304684 17428 485780 17456
rect 304684 17416 304690 17428
rect 485774 17416 485780 17428
rect 485832 17416 485838 17468
rect 304442 17348 304448 17400
rect 304500 17388 304506 17400
rect 485866 17388 485872 17400
rect 304500 17360 485872 17388
rect 304500 17348 304506 17360
rect 485866 17348 485872 17360
rect 485924 17348 485930 17400
rect 302050 17320 302056 17332
rect 302011 17292 302056 17320
rect 302050 17280 302056 17292
rect 302108 17280 302114 17332
rect 304534 17280 304540 17332
rect 304592 17320 304598 17332
rect 488534 17320 488540 17332
rect 304592 17292 488540 17320
rect 304592 17280 304598 17292
rect 488534 17280 488540 17292
rect 488592 17280 488598 17332
rect 301958 17252 301964 17264
rect 301919 17224 301964 17252
rect 301958 17212 301964 17224
rect 302016 17212 302022 17264
rect 302142 17252 302148 17264
rect 302103 17224 302148 17252
rect 302142 17212 302148 17224
rect 302200 17212 302206 17264
rect 304718 17212 304724 17264
rect 304776 17252 304782 17264
rect 489914 17252 489920 17264
rect 304776 17224 489920 17252
rect 304776 17212 304782 17224
rect 489914 17212 489920 17224
rect 489972 17212 489978 17264
rect 278406 17184 278412 17196
rect 278367 17156 278412 17184
rect 278406 17144 278412 17156
rect 278464 17144 278470 17196
rect 278590 17184 278596 17196
rect 278551 17156 278596 17184
rect 278590 17144 278596 17156
rect 278648 17144 278654 17196
rect 285030 17144 285036 17196
rect 285088 17184 285094 17196
rect 390554 17184 390560 17196
rect 285088 17156 390560 17184
rect 285088 17144 285094 17156
rect 390554 17144 390560 17156
rect 390612 17144 390618 17196
rect 278222 17116 278228 17128
rect 278183 17088 278228 17116
rect 278222 17076 278228 17088
rect 278280 17076 278286 17128
rect 278314 17076 278320 17128
rect 278372 17116 278378 17128
rect 278498 17116 278504 17128
rect 278372 17088 278417 17116
rect 278459 17088 278504 17116
rect 278372 17076 278378 17088
rect 278498 17076 278504 17088
rect 278556 17076 278562 17128
rect 278682 17116 278688 17128
rect 278643 17088 278688 17116
rect 278682 17076 278688 17088
rect 278740 17076 278746 17128
rect 283834 17076 283840 17128
rect 283892 17116 283898 17128
rect 387794 17116 387800 17128
rect 283892 17088 387800 17116
rect 283892 17076 283898 17088
rect 387794 17076 387800 17088
rect 387852 17076 387858 17128
rect 274082 17008 274088 17060
rect 274140 17048 274146 17060
rect 339770 17048 339776 17060
rect 274140 17020 339776 17048
rect 274140 17008 274146 17020
rect 339770 17008 339776 17020
rect 339828 17008 339834 17060
rect 274266 16940 274272 16992
rect 274324 16980 274330 16992
rect 339678 16980 339684 16992
rect 274324 16952 339684 16980
rect 274324 16940 274330 16952
rect 339678 16940 339684 16952
rect 339736 16940 339742 16992
rect 274174 16872 274180 16924
rect 274232 16912 274238 16924
rect 336734 16912 336740 16924
rect 274232 16884 336740 16912
rect 274232 16872 274238 16884
rect 336734 16872 336740 16884
rect 336792 16872 336798 16924
rect 505002 16872 505008 16924
rect 505060 16912 505066 16924
rect 511902 16912 511908 16924
rect 505060 16884 511908 16912
rect 505060 16872 505066 16884
rect 511902 16872 511908 16884
rect 511960 16872 511966 16924
rect 272794 16804 272800 16856
rect 272852 16844 272858 16856
rect 335354 16844 335360 16856
rect 272852 16816 335360 16844
rect 272852 16804 272858 16816
rect 335354 16804 335360 16816
rect 335412 16804 335418 16856
rect 272702 16736 272708 16788
rect 272760 16776 272766 16788
rect 332778 16776 332784 16788
rect 272760 16748 332784 16776
rect 272760 16736 272766 16748
rect 332778 16736 332784 16748
rect 332836 16736 332842 16788
rect 268746 16708 268752 16720
rect 268707 16680 268752 16708
rect 268746 16668 268752 16680
rect 268804 16668 268810 16720
rect 268930 16708 268936 16720
rect 268891 16680 268936 16708
rect 268930 16668 268936 16680
rect 268988 16668 268994 16720
rect 272886 16668 272892 16720
rect 272944 16708 272950 16720
rect 331306 16708 331312 16720
rect 272944 16680 331312 16708
rect 272944 16668 272950 16680
rect 331306 16668 331312 16680
rect 331364 16668 331370 16720
rect 394694 16668 394700 16720
rect 394752 16708 394758 16720
rect 404262 16708 404268 16720
rect 394752 16680 404268 16708
rect 394752 16668 394758 16680
rect 404262 16668 404268 16680
rect 404320 16668 404326 16720
rect 268838 16640 268844 16652
rect 268799 16612 268844 16640
rect 268838 16600 268844 16612
rect 268896 16600 268902 16652
rect 269022 16640 269028 16652
rect 268983 16612 269028 16640
rect 269022 16600 269028 16612
rect 269080 16600 269086 16652
rect 272978 16600 272984 16652
rect 273036 16640 273042 16652
rect 330110 16640 330116 16652
rect 273036 16612 330116 16640
rect 273036 16600 273042 16612
rect 330110 16600 330116 16612
rect 330168 16600 330174 16652
rect 330386 16600 330392 16652
rect 330444 16640 330450 16652
rect 330570 16640 330576 16652
rect 330444 16612 330576 16640
rect 330444 16600 330450 16612
rect 330570 16600 330576 16612
rect 330628 16600 330634 16652
rect 331858 16600 331864 16652
rect 331916 16640 331922 16652
rect 331950 16640 331956 16652
rect 331916 16612 331956 16640
rect 331916 16600 331922 16612
rect 331950 16600 331956 16612
rect 332008 16600 332014 16652
rect 437382 16600 437388 16652
rect 437440 16640 437446 16652
rect 442902 16640 442908 16652
rect 437440 16612 442908 16640
rect 437440 16600 437446 16612
rect 442902 16600 442908 16612
rect 442960 16600 442966 16652
rect 67542 16532 67548 16584
rect 67600 16572 67606 16584
rect 231121 16575 231179 16581
rect 231121 16572 231133 16575
rect 67600 16544 231133 16572
rect 67600 16532 67606 16544
rect 231121 16541 231133 16544
rect 231167 16541 231179 16575
rect 231121 16535 231179 16541
rect 231397 16575 231455 16581
rect 231397 16541 231409 16575
rect 231443 16572 231455 16575
rect 337010 16572 337016 16584
rect 231443 16544 337016 16572
rect 231443 16541 231455 16544
rect 231397 16535 231455 16541
rect 337010 16532 337016 16544
rect 337068 16532 337074 16584
rect 64782 16464 64788 16516
rect 64840 16504 64846 16516
rect 337102 16504 337108 16516
rect 64840 16476 337108 16504
rect 64840 16464 64846 16476
rect 337102 16464 337108 16476
rect 337160 16464 337166 16516
rect 60642 16396 60648 16448
rect 60700 16436 60706 16448
rect 335814 16436 335820 16448
rect 60700 16408 335820 16436
rect 60700 16396 60706 16408
rect 335814 16396 335820 16408
rect 335872 16396 335878 16448
rect 56502 16328 56508 16380
rect 56560 16368 56566 16380
rect 335538 16368 335544 16380
rect 56560 16340 335544 16368
rect 56560 16328 56566 16340
rect 335538 16328 335544 16340
rect 335596 16328 335602 16380
rect 53742 16260 53748 16312
rect 53800 16300 53806 16312
rect 334342 16300 334348 16312
rect 53800 16272 334348 16300
rect 53800 16260 53806 16272
rect 334342 16260 334348 16272
rect 334400 16260 334406 16312
rect 49602 16192 49608 16244
rect 49660 16232 49666 16244
rect 334066 16232 334072 16244
rect 49660 16204 334072 16232
rect 49660 16192 49666 16204
rect 334066 16192 334072 16204
rect 334124 16192 334130 16244
rect 345014 16192 345020 16244
rect 345072 16232 345078 16244
rect 346394 16232 346400 16244
rect 345072 16204 346400 16232
rect 345072 16192 345078 16204
rect 346394 16192 346400 16204
rect 346452 16192 346458 16244
rect 45462 16124 45468 16176
rect 45520 16164 45526 16176
rect 332870 16164 332876 16176
rect 45520 16136 332876 16164
rect 45520 16124 45526 16136
rect 332870 16124 332876 16136
rect 332928 16124 332934 16176
rect 41322 16056 41328 16108
rect 41380 16096 41386 16108
rect 331398 16096 331404 16108
rect 41380 16068 331404 16096
rect 41380 16056 41386 16068
rect 331398 16056 331404 16068
rect 331456 16056 331462 16108
rect 38562 15988 38568 16040
rect 38620 16028 38626 16040
rect 331490 16028 331496 16040
rect 38620 16000 331496 16028
rect 38620 15988 38626 16000
rect 331490 15988 331496 16000
rect 331548 15988 331554 16040
rect 34422 15920 34428 15972
rect 34480 15960 34486 15972
rect 330386 15960 330392 15972
rect 34480 15932 330392 15960
rect 34480 15920 34486 15932
rect 330386 15920 330392 15932
rect 330444 15920 330450 15972
rect 30282 15852 30288 15904
rect 30340 15892 30346 15904
rect 330202 15892 330208 15904
rect 30340 15864 330208 15892
rect 30340 15852 30346 15864
rect 330202 15852 330208 15864
rect 330260 15852 330266 15904
rect 95142 15784 95148 15836
rect 95200 15824 95206 15836
rect 342438 15824 342444 15836
rect 95200 15796 342444 15824
rect 95200 15784 95206 15796
rect 342438 15784 342444 15796
rect 342496 15784 342502 15836
rect 99190 15716 99196 15768
rect 99248 15756 99254 15768
rect 343726 15756 343732 15768
rect 99248 15728 343732 15756
rect 99248 15716 99254 15728
rect 343726 15716 343732 15728
rect 343784 15716 343790 15768
rect 102042 15648 102048 15700
rect 102100 15688 102106 15700
rect 344094 15688 344100 15700
rect 102100 15660 344100 15688
rect 102100 15648 102106 15660
rect 344094 15648 344100 15660
rect 344152 15648 344158 15700
rect 106182 15580 106188 15632
rect 106240 15620 106246 15632
rect 345106 15620 345112 15632
rect 106240 15592 345112 15620
rect 106240 15580 106246 15592
rect 345106 15580 345112 15592
rect 345164 15580 345170 15632
rect 108942 15512 108948 15564
rect 109000 15552 109006 15564
rect 345198 15552 345204 15564
rect 109000 15524 345204 15552
rect 109000 15512 109006 15524
rect 345198 15512 345204 15524
rect 345256 15512 345262 15564
rect 113082 15444 113088 15496
rect 113140 15484 113146 15496
rect 346946 15484 346952 15496
rect 113140 15456 346952 15484
rect 113140 15444 113146 15456
rect 346946 15444 346952 15456
rect 347004 15444 347010 15496
rect 117222 15376 117228 15428
rect 117280 15416 117286 15428
rect 348418 15416 348424 15428
rect 117280 15388 348424 15416
rect 117280 15376 117286 15388
rect 348418 15376 348424 15388
rect 348476 15376 348482 15428
rect 119982 15308 119988 15360
rect 120040 15348 120046 15360
rect 348050 15348 348056 15360
rect 120040 15320 348056 15348
rect 120040 15308 120046 15320
rect 348050 15308 348056 15320
rect 348108 15308 348114 15360
rect 124122 15240 124128 15292
rect 124180 15280 124186 15292
rect 349338 15280 349344 15292
rect 124180 15252 349344 15280
rect 124180 15240 124186 15252
rect 349338 15240 349344 15252
rect 349396 15240 349402 15292
rect 301958 15212 301964 15224
rect 301919 15184 301964 15212
rect 301958 15172 301964 15184
rect 302016 15172 302022 15224
rect 302142 15212 302148 15224
rect 302103 15184 302148 15212
rect 302142 15172 302148 15184
rect 302200 15172 302206 15224
rect 304626 15212 304632 15224
rect 304587 15184 304632 15212
rect 304626 15172 304632 15184
rect 304684 15172 304690 15224
rect 304902 15212 304908 15224
rect 304863 15184 304908 15212
rect 304902 15172 304908 15184
rect 304960 15172 304966 15224
rect 307202 15212 307208 15224
rect 307163 15184 307208 15212
rect 307202 15172 307208 15184
rect 307260 15172 307266 15224
rect 329098 15212 329104 15224
rect 329059 15184 329104 15212
rect 329098 15172 329104 15184
rect 329156 15172 329162 15224
rect 302050 15144 302056 15156
rect 302011 15116 302056 15144
rect 302050 15104 302056 15116
rect 302108 15104 302114 15156
rect 303154 15104 303160 15156
rect 303212 15144 303218 15156
rect 477494 15144 477500 15156
rect 303212 15116 477500 15144
rect 303212 15104 303218 15116
rect 477494 15104 477500 15116
rect 477552 15104 477558 15156
rect 303246 15036 303252 15088
rect 303304 15076 303310 15088
rect 481634 15076 481640 15088
rect 303304 15048 481640 15076
rect 303304 15036 303310 15048
rect 481634 15036 481640 15048
rect 481692 15036 481698 15088
rect 91002 14968 91008 15020
rect 91060 15008 91066 15020
rect 342898 15008 342904 15020
rect 91060 14980 342904 15008
rect 91060 14968 91066 14980
rect 342898 14968 342904 14980
rect 342956 14968 342962 15020
rect 88242 14900 88248 14952
rect 88300 14940 88306 14952
rect 340966 14940 340972 14952
rect 88300 14912 340972 14940
rect 88300 14900 88306 14912
rect 340966 14900 340972 14912
rect 341024 14900 341030 14952
rect 84102 14832 84108 14884
rect 84160 14872 84166 14884
rect 341242 14872 341248 14884
rect 84160 14844 341248 14872
rect 84160 14832 84166 14844
rect 341242 14832 341248 14844
rect 341300 14832 341306 14884
rect 81342 14764 81348 14816
rect 81400 14804 81406 14816
rect 339954 14804 339960 14816
rect 81400 14776 339960 14804
rect 81400 14764 81406 14776
rect 339954 14764 339960 14776
rect 340012 14764 340018 14816
rect 77202 14696 77208 14748
rect 77260 14736 77266 14748
rect 339586 14736 339592 14748
rect 77260 14708 339592 14736
rect 77260 14696 77266 14708
rect 339586 14696 339592 14708
rect 339644 14696 339650 14748
rect 73062 14628 73068 14680
rect 73120 14668 73126 14680
rect 338298 14668 338304 14680
rect 73120 14640 338304 14668
rect 73120 14628 73126 14640
rect 338298 14628 338304 14640
rect 338356 14628 338362 14680
rect 70302 14560 70308 14612
rect 70360 14600 70366 14612
rect 338206 14600 338212 14612
rect 70360 14572 338212 14600
rect 70360 14560 70366 14572
rect 338206 14560 338212 14572
rect 338264 14560 338270 14612
rect 66162 14492 66168 14544
rect 66220 14532 66226 14544
rect 336826 14532 336832 14544
rect 66220 14504 336832 14532
rect 66220 14492 66226 14504
rect 336826 14492 336832 14504
rect 336884 14492 336890 14544
rect 63402 14424 63408 14476
rect 63460 14464 63466 14476
rect 337286 14464 337292 14476
rect 63460 14436 337292 14464
rect 63460 14424 63466 14436
rect 337286 14424 337292 14436
rect 337344 14424 337350 14476
rect 301777 14399 301835 14405
rect 301777 14365 301789 14399
rect 301823 14396 301835 14399
rect 474734 14396 474740 14408
rect 301823 14368 474740 14396
rect 301823 14365 301835 14368
rect 301777 14359 301835 14365
rect 474734 14356 474740 14368
rect 474792 14356 474798 14408
rect 301869 14331 301927 14337
rect 301869 14297 301881 14331
rect 301915 14328 301927 14331
rect 470594 14328 470600 14340
rect 301915 14300 470600 14328
rect 301915 14297 301927 14300
rect 301869 14291 301927 14297
rect 470594 14288 470600 14300
rect 470652 14288 470658 14340
rect 300302 14220 300308 14272
rect 300360 14260 300366 14272
rect 467834 14260 467840 14272
rect 300360 14232 467840 14260
rect 300360 14220 300366 14232
rect 467834 14220 467840 14232
rect 467892 14220 467898 14272
rect 300394 14152 300400 14204
rect 300452 14192 300458 14204
rect 463694 14192 463700 14204
rect 300452 14164 463700 14192
rect 300452 14152 300458 14164
rect 463694 14152 463700 14164
rect 463752 14152 463758 14204
rect 299014 14084 299020 14136
rect 299072 14124 299078 14136
rect 459554 14124 459560 14136
rect 299072 14096 459560 14124
rect 299072 14084 299078 14096
rect 459554 14084 459560 14096
rect 459612 14084 459618 14136
rect 300673 14059 300731 14065
rect 300673 14025 300685 14059
rect 300719 14056 300731 14059
rect 456794 14056 456800 14068
rect 300719 14028 456800 14056
rect 300719 14025 300731 14028
rect 300673 14019 300731 14025
rect 456794 14016 456800 14028
rect 456852 14016 456858 14068
rect 297545 13991 297603 13997
rect 297545 13957 297557 13991
rect 297591 13988 297603 13991
rect 452654 13988 452660 14000
rect 297591 13960 452660 13988
rect 297591 13957 297603 13960
rect 297545 13951 297603 13957
rect 452654 13948 452660 13960
rect 452712 13948 452718 14000
rect 296162 13880 296168 13932
rect 296220 13920 296226 13932
rect 449894 13920 449900 13932
rect 296220 13892 449900 13920
rect 296220 13880 296226 13892
rect 449894 13880 449900 13892
rect 449952 13880 449958 13932
rect 296254 13812 296260 13864
rect 296312 13852 296318 13864
rect 445754 13852 445760 13864
rect 296312 13824 445760 13852
rect 296312 13812 296318 13824
rect 445754 13812 445760 13824
rect 445812 13812 445818 13864
rect 281074 13744 281080 13796
rect 281132 13784 281138 13796
rect 373994 13784 374000 13796
rect 281132 13756 374000 13784
rect 281132 13744 281138 13756
rect 373994 13744 374000 13756
rect 374052 13744 374058 13796
rect 283558 13676 283564 13728
rect 283616 13716 283622 13728
rect 378134 13716 378140 13728
rect 283616 13688 378140 13716
rect 283616 13676 283622 13688
rect 378134 13676 378140 13688
rect 378192 13676 378198 13728
rect 282454 13608 282460 13660
rect 282512 13648 282518 13660
rect 382274 13648 382280 13660
rect 282512 13620 382280 13648
rect 282512 13608 282518 13620
rect 382274 13608 382280 13620
rect 382332 13608 382338 13660
rect 283926 13540 283932 13592
rect 283984 13580 283990 13592
rect 385034 13580 385040 13592
rect 283984 13552 385040 13580
rect 283984 13540 283990 13552
rect 385034 13540 385040 13552
rect 385092 13540 385098 13592
rect 284018 13472 284024 13524
rect 284076 13512 284082 13524
rect 389174 13512 389180 13524
rect 284076 13484 389180 13512
rect 284076 13472 284082 13484
rect 389174 13472 389180 13484
rect 389232 13472 389238 13524
rect 285306 13404 285312 13456
rect 285364 13444 285370 13456
rect 391934 13444 391940 13456
rect 285364 13416 391940 13444
rect 285364 13404 285370 13416
rect 391934 13404 391940 13416
rect 391992 13404 391998 13456
rect 285214 13336 285220 13388
rect 285272 13376 285278 13388
rect 396074 13376 396080 13388
rect 285272 13348 396080 13376
rect 285272 13336 285278 13348
rect 396074 13336 396080 13348
rect 396132 13336 396138 13388
rect 286502 13268 286508 13320
rect 286560 13308 286566 13320
rect 400214 13308 400220 13320
rect 286560 13280 400220 13308
rect 286560 13268 286566 13280
rect 400214 13268 400220 13280
rect 400272 13268 400278 13320
rect 287974 13200 287980 13252
rect 288032 13240 288038 13252
rect 402974 13240 402980 13252
rect 288032 13212 402980 13240
rect 288032 13200 288038 13212
rect 402974 13200 402980 13212
rect 403032 13200 403038 13252
rect 268930 13172 268936 13184
rect 268891 13144 268936 13172
rect 268930 13132 268936 13144
rect 268988 13132 268994 13184
rect 287790 13132 287796 13184
rect 287848 13172 287854 13184
rect 407114 13172 407120 13184
rect 287848 13144 407120 13172
rect 287848 13132 287854 13144
rect 407114 13132 407120 13144
rect 407172 13132 407178 13184
rect 268746 13104 268752 13116
rect 268707 13076 268752 13104
rect 268746 13064 268752 13076
rect 268804 13064 268810 13116
rect 269022 13104 269028 13116
rect 268983 13076 269028 13104
rect 269022 13064 269028 13076
rect 269080 13064 269086 13116
rect 278682 13104 278688 13116
rect 278643 13076 278688 13104
rect 278682 13064 278688 13076
rect 278740 13064 278746 13116
rect 289170 13064 289176 13116
rect 289228 13104 289234 13116
rect 409874 13104 409880 13116
rect 289228 13076 409880 13104
rect 289228 13064 289234 13076
rect 409874 13064 409880 13076
rect 409932 13064 409938 13116
rect 280982 12996 280988 13048
rect 281040 13036 281046 13048
rect 371234 13036 371240 13048
rect 281040 13008 371240 13036
rect 281040 12996 281046 13008
rect 371234 12996 371240 13008
rect 371292 12996 371298 13048
rect 279694 12928 279700 12980
rect 279752 12968 279758 12980
rect 367094 12968 367100 12980
rect 279752 12940 367100 12968
rect 279752 12928 279758 12940
rect 367094 12928 367100 12940
rect 367152 12928 367158 12980
rect 279786 12860 279792 12912
rect 279844 12900 279850 12912
rect 364334 12900 364340 12912
rect 279844 12872 364340 12900
rect 279844 12860 279850 12872
rect 364334 12860 364340 12872
rect 364392 12860 364398 12912
rect 278317 12835 278375 12841
rect 278317 12801 278329 12835
rect 278363 12832 278375 12835
rect 360194 12832 360200 12844
rect 278363 12804 360200 12832
rect 278363 12801 278375 12804
rect 278317 12795 278375 12801
rect 360194 12792 360200 12804
rect 360252 12792 360258 12844
rect 278225 12767 278283 12773
rect 278225 12733 278237 12767
rect 278271 12764 278283 12767
rect 356054 12764 356060 12776
rect 278271 12736 356060 12764
rect 278271 12733 278283 12736
rect 278225 12727 278283 12733
rect 356054 12724 356060 12736
rect 356112 12724 356118 12776
rect 276934 12656 276940 12708
rect 276992 12696 276998 12708
rect 353294 12696 353300 12708
rect 276992 12668 353300 12696
rect 276992 12656 276998 12668
rect 353294 12656 353300 12668
rect 353352 12656 353358 12708
rect 276842 12588 276848 12640
rect 276900 12628 276906 12640
rect 349154 12628 349160 12640
rect 276900 12600 349160 12628
rect 276900 12588 276906 12600
rect 349154 12588 349160 12600
rect 349212 12588 349218 12640
rect 268838 12560 268844 12572
rect 268799 12532 268844 12560
rect 268838 12520 268844 12532
rect 268896 12520 268902 12572
rect 275554 12520 275560 12572
rect 275612 12560 275618 12572
rect 346578 12560 346584 12572
rect 275612 12532 346584 12560
rect 275612 12520 275618 12532
rect 346578 12520 346584 12532
rect 346636 12520 346642 12572
rect 244458 12492 244464 12504
rect 244384 12464 244464 12492
rect 244384 12436 244412 12464
rect 244458 12452 244464 12464
rect 244516 12452 244522 12504
rect 244918 12492 244924 12504
rect 244844 12464 244924 12492
rect 244844 12436 244872 12464
rect 244918 12452 244924 12464
rect 244976 12452 244982 12504
rect 274358 12452 274364 12504
rect 274416 12492 274422 12504
rect 342622 12492 342628 12504
rect 274416 12464 342628 12492
rect 274416 12452 274422 12464
rect 342622 12452 342628 12464
rect 342680 12452 342686 12504
rect 244366 12384 244372 12436
rect 244424 12384 244430 12436
rect 244826 12384 244832 12436
rect 244884 12384 244890 12436
rect 275554 12384 275560 12436
rect 275612 12424 275618 12436
rect 275830 12424 275836 12436
rect 275612 12396 275836 12424
rect 275612 12384 275618 12396
rect 275830 12384 275836 12396
rect 275888 12384 275894 12436
rect 307018 12384 307024 12436
rect 307076 12424 307082 12436
rect 307294 12424 307300 12436
rect 307076 12396 307300 12424
rect 307076 12384 307082 12396
rect 307294 12384 307300 12396
rect 307352 12384 307358 12436
rect 308490 12384 308496 12436
rect 308548 12424 308554 12436
rect 308582 12424 308588 12436
rect 308548 12396 308588 12424
rect 308548 12384 308554 12396
rect 308582 12384 308588 12396
rect 308640 12384 308646 12436
rect 309962 12384 309968 12436
rect 310020 12424 310026 12436
rect 310054 12424 310060 12436
rect 310020 12396 310060 12424
rect 310020 12384 310026 12396
rect 310054 12384 310060 12396
rect 310112 12384 310118 12436
rect 520274 12424 520280 12436
rect 311360 12396 520280 12424
rect 311360 12368 311388 12396
rect 520274 12384 520280 12396
rect 520332 12384 520338 12436
rect 311342 12316 311348 12368
rect 311400 12316 311406 12368
rect 312722 12316 312728 12368
rect 312780 12356 312786 12368
rect 524414 12356 524420 12368
rect 312780 12328 524420 12356
rect 312780 12316 312786 12328
rect 524414 12316 524420 12328
rect 524472 12316 524478 12368
rect 312814 12248 312820 12300
rect 312872 12288 312878 12300
rect 528554 12288 528560 12300
rect 312872 12260 528560 12288
rect 312872 12248 312878 12260
rect 528554 12248 528560 12260
rect 528612 12248 528618 12300
rect 314378 12180 314384 12232
rect 314436 12220 314442 12232
rect 531314 12220 531320 12232
rect 314436 12192 531320 12220
rect 314436 12180 314442 12192
rect 531314 12180 531320 12192
rect 531372 12180 531378 12232
rect 314286 12112 314292 12164
rect 314344 12152 314350 12164
rect 535454 12152 535460 12164
rect 314344 12124 535460 12152
rect 314344 12112 314350 12124
rect 535454 12112 535460 12124
rect 535512 12112 535518 12164
rect 278590 12084 278596 12096
rect 278551 12056 278596 12084
rect 278590 12044 278596 12056
rect 278648 12044 278654 12096
rect 315666 12044 315672 12096
rect 315724 12084 315730 12096
rect 538214 12084 538220 12096
rect 315724 12056 538220 12084
rect 315724 12044 315730 12056
rect 538214 12044 538220 12056
rect 538272 12044 538278 12096
rect 315758 11976 315764 12028
rect 315816 12016 315822 12028
rect 542354 12016 542360 12028
rect 315816 11988 542360 12016
rect 315816 11976 315822 11988
rect 542354 11976 542360 11988
rect 542412 11976 542418 12028
rect 317046 11908 317052 11960
rect 317104 11948 317110 11960
rect 546494 11948 546500 11960
rect 317104 11920 546500 11948
rect 317104 11908 317110 11920
rect 546494 11908 546500 11920
rect 546552 11908 546558 11960
rect 316862 11840 316868 11892
rect 316920 11880 316926 11892
rect 549254 11880 549260 11892
rect 316920 11852 549260 11880
rect 316920 11840 316926 11852
rect 549254 11840 549260 11852
rect 549312 11840 549318 11892
rect 318150 11772 318156 11824
rect 318208 11812 318214 11824
rect 553394 11812 553400 11824
rect 318208 11784 553400 11812
rect 318208 11772 318214 11784
rect 553394 11772 553400 11784
rect 553452 11772 553458 11824
rect 318334 11704 318340 11756
rect 318392 11744 318398 11756
rect 556154 11744 556160 11756
rect 318392 11716 556160 11744
rect 318392 11704 318398 11716
rect 556154 11704 556160 11716
rect 556212 11704 556218 11756
rect 311434 11636 311440 11688
rect 311492 11676 311498 11688
rect 517514 11676 517520 11688
rect 311492 11648 517520 11676
rect 311492 11636 311498 11648
rect 517514 11636 517520 11648
rect 517572 11636 517578 11688
rect 309962 11568 309968 11620
rect 310020 11608 310026 11620
rect 513374 11608 513380 11620
rect 310020 11580 513380 11608
rect 310020 11568 310026 11580
rect 513374 11568 513380 11580
rect 513432 11568 513438 11620
rect 308674 11500 308680 11552
rect 308732 11540 308738 11552
rect 510614 11540 510620 11552
rect 308732 11512 510620 11540
rect 308732 11500 308738 11512
rect 510614 11500 510620 11512
rect 510672 11500 510678 11552
rect 308490 11432 308496 11484
rect 308548 11472 308554 11484
rect 506474 11472 506480 11484
rect 308548 11444 506480 11472
rect 308548 11432 308554 11444
rect 506474 11432 506480 11444
rect 506532 11432 506538 11484
rect 307205 11407 307263 11413
rect 307205 11373 307217 11407
rect 307251 11404 307263 11407
rect 502334 11404 502340 11416
rect 307251 11376 502340 11404
rect 307251 11373 307263 11376
rect 307205 11367 307263 11373
rect 502334 11364 502340 11376
rect 502392 11364 502398 11416
rect 307018 11296 307024 11348
rect 307076 11336 307082 11348
rect 499574 11336 499580 11348
rect 307076 11308 499580 11336
rect 307076 11296 307082 11308
rect 499574 11296 499580 11308
rect 499632 11296 499638 11348
rect 306006 11228 306012 11280
rect 306064 11268 306070 11280
rect 495434 11268 495440 11280
rect 306064 11240 495440 11268
rect 306064 11228 306070 11240
rect 495434 11228 495440 11240
rect 495492 11228 495498 11280
rect 271506 11160 271512 11212
rect 271564 11200 271570 11212
rect 328822 11200 328828 11212
rect 271564 11172 328828 11200
rect 271564 11160 271570 11172
rect 328822 11160 328828 11172
rect 328880 11160 328886 11212
rect 271414 11092 271420 11144
rect 271472 11132 271478 11144
rect 324406 11132 324412 11144
rect 271472 11104 324412 11132
rect 271472 11092 271478 11104
rect 324406 11092 324412 11104
rect 324464 11092 324470 11144
rect 314378 11024 314384 11076
rect 314436 11064 314442 11076
rect 314562 11064 314568 11076
rect 314436 11036 314568 11064
rect 314436 11024 314442 11036
rect 314562 11024 314568 11036
rect 314620 11024 314626 11076
rect 322474 11024 322480 11076
rect 322532 11064 322538 11076
rect 322658 11064 322664 11076
rect 322532 11036 322664 11064
rect 322532 11024 322538 11036
rect 322658 11024 322664 11036
rect 322716 11024 322722 11076
rect 345382 11064 345388 11076
rect 345343 11036 345388 11064
rect 345382 11024 345388 11036
rect 345440 11024 345446 11076
rect 292206 10956 292212 11008
rect 292264 10996 292270 11008
rect 426434 10996 426440 11008
rect 292264 10968 426440 10996
rect 292264 10956 292270 10968
rect 426434 10956 426440 10968
rect 426492 10956 426498 11008
rect 293862 10888 293868 10940
rect 293920 10928 293926 10940
rect 430574 10928 430580 10940
rect 293920 10900 430580 10928
rect 293920 10888 293926 10900
rect 430574 10888 430580 10900
rect 430632 10888 430638 10940
rect 293770 10820 293776 10872
rect 293828 10860 293834 10872
rect 433426 10860 433432 10872
rect 293828 10832 433432 10860
rect 293828 10820 293834 10832
rect 433426 10820 433432 10832
rect 433484 10820 433490 10872
rect 295242 10752 295248 10804
rect 295300 10792 295306 10804
rect 437474 10792 437480 10804
rect 295300 10764 437480 10792
rect 295300 10752 295306 10764
rect 437474 10752 437480 10764
rect 437532 10752 437538 10804
rect 295150 10684 295156 10736
rect 295208 10724 295214 10736
rect 441614 10724 441620 10736
rect 295208 10696 441620 10724
rect 295208 10684 295214 10696
rect 441614 10684 441620 10696
rect 441672 10684 441678 10736
rect 296346 10616 296352 10668
rect 296404 10656 296410 10668
rect 444374 10656 444380 10668
rect 296404 10628 444380 10656
rect 296404 10616 296410 10628
rect 444374 10616 444380 10628
rect 444432 10616 444438 10668
rect 296438 10548 296444 10600
rect 296496 10588 296502 10600
rect 448514 10588 448520 10600
rect 296496 10560 448520 10588
rect 296496 10548 296502 10560
rect 448514 10548 448520 10560
rect 448572 10548 448578 10600
rect 297726 10480 297732 10532
rect 297784 10520 297790 10532
rect 451274 10520 451280 10532
rect 297784 10492 451280 10520
rect 297784 10480 297790 10492
rect 451274 10480 451280 10492
rect 451332 10480 451338 10532
rect 297818 10412 297824 10464
rect 297876 10452 297882 10464
rect 455414 10452 455420 10464
rect 297876 10424 455420 10452
rect 297876 10412 297882 10424
rect 455414 10412 455420 10424
rect 455472 10412 455478 10464
rect 299198 10344 299204 10396
rect 299256 10384 299262 10396
rect 459646 10384 459652 10396
rect 299256 10356 459652 10384
rect 299256 10344 299262 10356
rect 459646 10344 459652 10356
rect 459704 10344 459710 10396
rect 299106 10276 299112 10328
rect 299164 10316 299170 10328
rect 462314 10316 462320 10328
rect 299164 10288 462320 10316
rect 299164 10276 299170 10288
rect 462314 10276 462320 10288
rect 462372 10276 462378 10328
rect 292298 10208 292304 10260
rect 292356 10248 292362 10260
rect 423674 10248 423680 10260
rect 292356 10220 423680 10248
rect 292356 10208 292362 10220
rect 423674 10208 423680 10220
rect 423732 10208 423738 10260
rect 290918 10140 290924 10192
rect 290976 10180 290982 10192
rect 419534 10180 419540 10192
rect 290976 10152 419540 10180
rect 290976 10140 290982 10152
rect 419534 10140 419540 10152
rect 419592 10140 419598 10192
rect 289446 10072 289452 10124
rect 289504 10112 289510 10124
rect 416866 10112 416872 10124
rect 289504 10084 416872 10112
rect 289504 10072 289510 10084
rect 416866 10072 416872 10084
rect 416924 10072 416930 10124
rect 289538 10004 289544 10056
rect 289596 10044 289602 10056
rect 412634 10044 412640 10056
rect 289596 10016 412640 10044
rect 289596 10004 289602 10016
rect 412634 10004 412640 10016
rect 412692 10004 412698 10056
rect 288158 9936 288164 9988
rect 288216 9976 288222 9988
rect 408494 9976 408500 9988
rect 288216 9948 408500 9976
rect 288216 9936 288222 9948
rect 408494 9936 408500 9948
rect 408552 9936 408558 9988
rect 288066 9868 288072 9920
rect 288124 9908 288130 9920
rect 405734 9908 405740 9920
rect 288124 9880 405740 9908
rect 288124 9868 288130 9880
rect 405734 9868 405740 9880
rect 405792 9868 405798 9920
rect 288434 9800 288440 9852
rect 288492 9840 288498 9852
rect 401594 9840 401600 9852
rect 288492 9812 401600 9840
rect 288492 9800 288498 9812
rect 401594 9800 401600 9812
rect 401652 9800 401658 9852
rect 286778 9732 286784 9784
rect 286836 9772 286842 9784
rect 398834 9772 398840 9784
rect 286836 9744 398840 9772
rect 286836 9732 286842 9744
rect 398834 9732 398840 9744
rect 398892 9732 398898 9784
rect 107473 9707 107531 9713
rect 107473 9673 107485 9707
rect 107519 9704 107531 9707
rect 107746 9704 107752 9716
rect 107519 9676 107752 9704
rect 107519 9673 107531 9676
rect 107473 9667 107531 9673
rect 107746 9664 107752 9676
rect 107804 9664 107810 9716
rect 232590 9664 232596 9716
rect 232648 9704 232654 9716
rect 232774 9704 232780 9716
rect 232648 9676 232780 9704
rect 232648 9664 232654 9676
rect 232774 9664 232780 9676
rect 232832 9664 232838 9716
rect 267090 9664 267096 9716
rect 267148 9704 267154 9716
rect 267182 9704 267188 9716
rect 267148 9676 267188 9704
rect 267148 9664 267154 9676
rect 267182 9664 267188 9676
rect 267240 9664 267246 9716
rect 268562 9664 268568 9716
rect 268620 9704 268626 9716
rect 268654 9704 268660 9716
rect 268620 9676 268660 9704
rect 268620 9664 268626 9676
rect 268654 9664 268660 9676
rect 268712 9664 268718 9716
rect 285398 9664 285404 9716
rect 285456 9704 285462 9716
rect 394694 9704 394700 9716
rect 285456 9676 394700 9704
rect 285456 9664 285462 9676
rect 394694 9664 394700 9676
rect 394752 9664 394758 9716
rect 90913 9639 90971 9645
rect 90913 9605 90925 9639
rect 90959 9636 90971 9639
rect 91002 9636 91008 9648
rect 90959 9608 91008 9636
rect 90959 9605 90971 9608
rect 90913 9599 90971 9605
rect 91002 9596 91008 9608
rect 91060 9596 91066 9648
rect 100481 9639 100539 9645
rect 100481 9605 100493 9639
rect 100527 9636 100539 9639
rect 100662 9636 100668 9648
rect 100527 9608 100668 9636
rect 100527 9605 100539 9608
rect 100481 9599 100539 9605
rect 100662 9596 100668 9608
rect 100720 9596 100726 9648
rect 108761 9639 108819 9645
rect 108761 9605 108773 9639
rect 108807 9636 108819 9639
rect 108942 9636 108948 9648
rect 108807 9608 108948 9636
rect 108807 9605 108819 9608
rect 108761 9599 108819 9605
rect 108942 9596 108948 9608
rect 109000 9596 109006 9648
rect 278409 9639 278467 9645
rect 278409 9605 278421 9639
rect 278455 9636 278467 9639
rect 359734 9636 359740 9648
rect 278455 9608 359740 9636
rect 278455 9605 278467 9608
rect 278409 9599 278467 9605
rect 359734 9596 359740 9608
rect 359792 9596 359798 9648
rect 278501 9571 278559 9577
rect 278501 9537 278513 9571
rect 278547 9568 278559 9571
rect 363322 9568 363328 9580
rect 278547 9540 363328 9568
rect 278547 9537 278559 9540
rect 278501 9531 278559 9537
rect 363322 9528 363328 9540
rect 363380 9528 363386 9580
rect 167086 9460 167092 9512
rect 167144 9500 167150 9512
rect 237926 9500 237932 9512
rect 167144 9472 237932 9500
rect 167144 9460 167150 9472
rect 237926 9460 237932 9472
rect 237984 9460 237990 9512
rect 279878 9460 279884 9512
rect 279936 9500 279942 9512
rect 366910 9500 366916 9512
rect 279936 9472 366916 9500
rect 279936 9460 279942 9472
rect 366910 9460 366916 9472
rect 366968 9460 366974 9512
rect 169386 9392 169392 9444
rect 169444 9432 169450 9444
rect 239214 9432 239220 9444
rect 169444 9404 239220 9432
rect 169444 9392 169450 9404
rect 239214 9392 239220 9404
rect 239272 9392 239278 9444
rect 281258 9392 281264 9444
rect 281316 9432 281322 9444
rect 370406 9432 370412 9444
rect 281316 9404 370412 9432
rect 281316 9392 281322 9404
rect 370406 9392 370412 9404
rect 370464 9392 370470 9444
rect 165890 9324 165896 9376
rect 165948 9364 165954 9376
rect 237466 9364 237472 9376
rect 165948 9336 237472 9364
rect 165948 9324 165954 9336
rect 237466 9324 237472 9336
rect 237524 9324 237530 9376
rect 281166 9324 281172 9376
rect 281224 9364 281230 9376
rect 374086 9364 374092 9376
rect 281224 9336 374092 9364
rect 281224 9324 281230 9336
rect 374086 9324 374092 9336
rect 374144 9324 374150 9376
rect 164694 9256 164700 9308
rect 164752 9296 164758 9308
rect 237742 9296 237748 9308
rect 164752 9268 237748 9296
rect 164752 9256 164758 9268
rect 237742 9256 237748 9268
rect 237800 9256 237806 9308
rect 282546 9256 282552 9308
rect 282604 9296 282610 9308
rect 377582 9296 377588 9308
rect 282604 9268 377588 9296
rect 282604 9256 282610 9268
rect 377582 9256 377588 9268
rect 377640 9256 377646 9308
rect 163498 9188 163504 9240
rect 163556 9228 163562 9240
rect 237650 9228 237656 9240
rect 163556 9200 237656 9228
rect 163556 9188 163562 9200
rect 237650 9188 237656 9200
rect 237708 9188 237714 9240
rect 282638 9188 282644 9240
rect 282696 9228 282702 9240
rect 381170 9228 381176 9240
rect 282696 9200 381176 9228
rect 282696 9188 282702 9200
rect 381170 9188 381176 9200
rect 381228 9188 381234 9240
rect 162302 9120 162308 9172
rect 162360 9160 162366 9172
rect 236638 9160 236644 9172
rect 162360 9132 236644 9160
rect 162360 9120 162366 9132
rect 236638 9120 236644 9132
rect 236696 9120 236702 9172
rect 268654 9120 268660 9172
rect 268712 9160 268718 9172
rect 314562 9160 314568 9172
rect 268712 9132 314568 9160
rect 268712 9120 268718 9132
rect 314562 9120 314568 9132
rect 314620 9120 314626 9172
rect 318058 9160 318064 9172
rect 314948 9132 318064 9160
rect 161106 9052 161112 9104
rect 161164 9092 161170 9104
rect 236454 9092 236460 9104
rect 161164 9064 236460 9092
rect 161164 9052 161170 9064
rect 236454 9052 236460 9064
rect 236512 9052 236518 9104
rect 270034 9052 270040 9104
rect 270092 9092 270098 9104
rect 314948 9092 314976 9132
rect 318058 9120 318064 9132
rect 318116 9120 318122 9172
rect 318518 9120 318524 9172
rect 318576 9160 318582 9172
rect 323121 9163 323179 9169
rect 318576 9132 322796 9160
rect 318576 9120 318582 9132
rect 270092 9064 314976 9092
rect 270092 9052 270098 9064
rect 317230 9052 317236 9104
rect 317288 9092 317294 9104
rect 322661 9095 322719 9101
rect 322661 9092 322673 9095
rect 317288 9064 322673 9092
rect 317288 9052 317294 9064
rect 322661 9061 322673 9064
rect 322707 9061 322719 9095
rect 322768 9092 322796 9132
rect 323121 9129 323133 9163
rect 323167 9160 323179 9163
rect 545298 9160 545304 9172
rect 323167 9132 545304 9160
rect 323167 9129 323179 9132
rect 323121 9123 323179 9129
rect 545298 9120 545304 9132
rect 545356 9120 545362 9172
rect 323029 9095 323087 9101
rect 322768 9064 322888 9092
rect 322661 9055 322719 9061
rect 128998 8984 129004 9036
rect 129056 9024 129062 9036
rect 230474 9024 230480 9036
rect 129056 8996 230480 9024
rect 129056 8984 129062 8996
rect 230474 8984 230480 8996
rect 230532 8984 230538 9036
rect 271598 8984 271604 9036
rect 271656 9024 271662 9036
rect 322753 9027 322811 9033
rect 322753 9024 322765 9027
rect 271656 8996 322765 9024
rect 271656 8984 271662 8996
rect 322753 8993 322765 8996
rect 322799 8993 322811 9027
rect 322860 9024 322888 9064
rect 323029 9061 323041 9095
rect 323075 9092 323087 9095
rect 324038 9092 324044 9104
rect 323075 9064 324044 9092
rect 323075 9061 323087 9064
rect 323029 9055 323087 9061
rect 324038 9052 324044 9064
rect 324096 9052 324102 9104
rect 552382 9092 552388 9104
rect 324148 9064 552388 9092
rect 324148 9024 324176 9064
rect 552382 9052 552388 9064
rect 552440 9052 552446 9104
rect 322860 8996 324176 9024
rect 324501 9027 324559 9033
rect 322753 8987 322811 8993
rect 324501 8993 324513 9027
rect 324547 9024 324559 9027
rect 577406 9024 577412 9036
rect 324547 8996 577412 9024
rect 324547 8993 324559 8996
rect 324501 8987 324559 8993
rect 577406 8984 577412 8996
rect 577464 8984 577470 9036
rect 126606 8916 126612 8968
rect 126664 8956 126670 8968
rect 229278 8956 229284 8968
rect 126664 8928 229284 8956
rect 126664 8916 126670 8928
rect 229278 8916 229284 8928
rect 229336 8916 229342 8968
rect 269942 8916 269948 8968
rect 270000 8956 270006 8968
rect 321646 8956 321652 8968
rect 270000 8928 321652 8956
rect 270000 8916 270006 8928
rect 321646 8916 321652 8928
rect 321704 8916 321710 8968
rect 322566 8916 322572 8968
rect 322624 8956 322630 8968
rect 324041 8959 324099 8965
rect 324041 8956 324053 8959
rect 322624 8928 324053 8956
rect 322624 8916 322630 8928
rect 324041 8925 324053 8928
rect 324087 8925 324099 8959
rect 324041 8919 324099 8925
rect 324130 8916 324136 8968
rect 324188 8956 324194 8968
rect 581086 8956 581092 8968
rect 324188 8928 581092 8956
rect 324188 8916 324194 8928
rect 581086 8916 581092 8928
rect 581144 8916 581150 8968
rect 277118 8848 277124 8900
rect 277176 8888 277182 8900
rect 356146 8888 356152 8900
rect 277176 8860 356152 8888
rect 277176 8848 277182 8860
rect 356146 8848 356152 8860
rect 356204 8848 356210 8900
rect 277026 8780 277032 8832
rect 277084 8820 277090 8832
rect 352558 8820 352564 8832
rect 277084 8792 352564 8820
rect 277084 8780 277090 8792
rect 352558 8780 352564 8792
rect 352616 8780 352622 8832
rect 275738 8712 275744 8764
rect 275796 8752 275802 8764
rect 349062 8752 349068 8764
rect 275796 8724 349068 8752
rect 275796 8712 275802 8724
rect 349062 8712 349068 8724
rect 349120 8712 349126 8764
rect 275646 8644 275652 8696
rect 275704 8684 275710 8696
rect 345474 8684 345480 8696
rect 275704 8656 345480 8684
rect 275704 8644 275710 8656
rect 345474 8644 345480 8656
rect 345532 8644 345538 8696
rect 274450 8576 274456 8628
rect 274508 8616 274514 8628
rect 341886 8616 341892 8628
rect 274508 8588 341892 8616
rect 274508 8576 274514 8588
rect 341886 8576 341892 8588
rect 341944 8576 341950 8628
rect 274542 8508 274548 8560
rect 274600 8548 274606 8560
rect 338298 8548 338304 8560
rect 274600 8520 338304 8548
rect 274600 8508 274606 8520
rect 338298 8508 338304 8520
rect 338356 8508 338362 8560
rect 273070 8440 273076 8492
rect 273128 8480 273134 8492
rect 334710 8480 334716 8492
rect 273128 8452 334716 8480
rect 273128 8440 273134 8452
rect 334710 8440 334716 8452
rect 334768 8440 334774 8492
rect 273162 8372 273168 8424
rect 273220 8412 273226 8424
rect 331214 8412 331220 8424
rect 273220 8384 331220 8412
rect 273220 8372 273226 8384
rect 331214 8372 331220 8384
rect 331272 8372 331278 8424
rect 271690 8304 271696 8356
rect 271748 8344 271754 8356
rect 327626 8344 327632 8356
rect 271748 8316 327632 8344
rect 271748 8304 271754 8316
rect 327626 8304 327632 8316
rect 327684 8304 327690 8356
rect 328454 8304 328460 8356
rect 328512 8344 328518 8356
rect 328914 8344 328920 8356
rect 328512 8316 328920 8344
rect 328512 8304 328518 8316
rect 328914 8304 328920 8316
rect 328972 8304 328978 8356
rect 345382 8344 345388 8356
rect 345343 8316 345388 8344
rect 345382 8304 345388 8316
rect 345440 8304 345446 8356
rect 196802 8236 196808 8288
rect 196860 8276 196866 8288
rect 244550 8276 244556 8288
rect 196860 8248 244556 8276
rect 196860 8236 196866 8248
rect 244550 8236 244556 8248
rect 244608 8236 244614 8288
rect 252922 8276 252928 8288
rect 252883 8248 252928 8276
rect 252922 8236 252928 8248
rect 252980 8236 252986 8288
rect 302142 8236 302148 8288
rect 302200 8276 302206 8288
rect 472710 8276 472716 8288
rect 302200 8248 472716 8276
rect 302200 8236 302206 8248
rect 472710 8236 472716 8248
rect 472768 8236 472774 8288
rect 193214 8168 193220 8220
rect 193272 8208 193278 8220
rect 243354 8208 243360 8220
rect 193272 8180 243360 8208
rect 193272 8168 193278 8180
rect 243354 8168 243360 8180
rect 243412 8168 243418 8220
rect 302050 8168 302056 8220
rect 302108 8208 302114 8220
rect 476298 8208 476304 8220
rect 302108 8180 476304 8208
rect 302108 8168 302114 8180
rect 476298 8168 476304 8180
rect 476356 8168 476362 8220
rect 189626 8100 189632 8152
rect 189684 8140 189690 8152
rect 243262 8140 243268 8152
rect 189684 8112 243268 8140
rect 189684 8100 189690 8112
rect 243262 8100 243268 8112
rect 243320 8100 243326 8152
rect 303522 8100 303528 8152
rect 303580 8140 303586 8152
rect 479886 8140 479892 8152
rect 303580 8112 479892 8140
rect 303580 8100 303586 8112
rect 479886 8100 479892 8112
rect 479944 8100 479950 8152
rect 186038 8032 186044 8084
rect 186096 8072 186102 8084
rect 241882 8072 241888 8084
rect 186096 8044 241888 8072
rect 186096 8032 186102 8044
rect 241882 8032 241888 8044
rect 241940 8032 241946 8084
rect 304902 8032 304908 8084
rect 304960 8072 304966 8084
rect 484578 8072 484584 8084
rect 304960 8044 484584 8072
rect 304960 8032 304966 8044
rect 484578 8032 484584 8044
rect 484636 8032 484642 8084
rect 182542 7964 182548 8016
rect 182600 8004 182606 8016
rect 241514 8004 241520 8016
rect 182600 7976 241520 8004
rect 182600 7964 182606 7976
rect 241514 7964 241520 7976
rect 241572 7964 241578 8016
rect 304810 7964 304816 8016
rect 304868 8004 304874 8016
rect 488166 8004 488172 8016
rect 304868 7976 488172 8004
rect 304868 7964 304874 7976
rect 488166 7964 488172 7976
rect 488224 7964 488230 8016
rect 178954 7896 178960 7948
rect 179012 7936 179018 7948
rect 240686 7936 240692 7948
rect 179012 7908 240692 7936
rect 179012 7896 179018 7908
rect 240686 7896 240692 7908
rect 240744 7896 240750 7948
rect 264514 7896 264520 7948
rect 264572 7936 264578 7948
rect 293126 7936 293132 7948
rect 264572 7908 293132 7936
rect 264572 7896 264578 7908
rect 293126 7896 293132 7908
rect 293184 7896 293190 7948
rect 306098 7896 306104 7948
rect 306156 7936 306162 7948
rect 491754 7936 491760 7948
rect 306156 7908 491760 7936
rect 306156 7896 306162 7908
rect 491754 7896 491760 7908
rect 491812 7896 491818 7948
rect 175366 7828 175372 7880
rect 175424 7868 175430 7880
rect 239122 7868 239128 7880
rect 175424 7840 239128 7868
rect 175424 7828 175430 7840
rect 239122 7828 239128 7840
rect 239180 7828 239186 7880
rect 265894 7828 265900 7880
rect 265952 7868 265958 7880
rect 296714 7868 296720 7880
rect 265952 7840 296720 7868
rect 265952 7828 265958 7840
rect 296714 7828 296720 7840
rect 296772 7828 296778 7880
rect 306190 7828 306196 7880
rect 306248 7868 306254 7880
rect 495342 7868 495348 7880
rect 306248 7840 495348 7868
rect 306248 7828 306254 7840
rect 495342 7828 495348 7840
rect 495400 7828 495406 7880
rect 171778 7760 171784 7812
rect 171836 7800 171842 7812
rect 239306 7800 239312 7812
rect 171836 7772 239312 7800
rect 171836 7760 171842 7772
rect 239306 7760 239312 7772
rect 239364 7760 239370 7812
rect 265802 7760 265808 7812
rect 265860 7800 265866 7812
rect 300302 7800 300308 7812
rect 265860 7772 300308 7800
rect 265860 7760 265866 7772
rect 300302 7760 300308 7772
rect 300360 7760 300366 7812
rect 307386 7760 307392 7812
rect 307444 7760 307450 7812
rect 307478 7760 307484 7812
rect 307536 7800 307542 7812
rect 498930 7800 498936 7812
rect 307536 7772 498936 7800
rect 307536 7760 307542 7772
rect 498930 7760 498936 7772
rect 498988 7760 498994 7812
rect 168190 7692 168196 7744
rect 168248 7732 168254 7744
rect 237374 7732 237380 7744
rect 168248 7704 237380 7732
rect 168248 7692 168254 7704
rect 237374 7692 237380 7704
rect 237432 7692 237438 7744
rect 267182 7692 267188 7744
rect 267240 7732 267246 7744
rect 303798 7732 303804 7744
rect 267240 7704 303804 7732
rect 267240 7692 267246 7704
rect 303798 7692 303804 7704
rect 303856 7692 303862 7744
rect 307404 7732 307432 7760
rect 502426 7732 502432 7744
rect 307404 7704 502432 7732
rect 502426 7692 502432 7704
rect 502484 7692 502490 7744
rect 157518 7624 157524 7676
rect 157576 7664 157582 7676
rect 236270 7664 236276 7676
rect 157576 7636 236276 7664
rect 157576 7624 157582 7636
rect 236270 7624 236276 7636
rect 236328 7624 236334 7676
rect 267274 7624 267280 7676
rect 267332 7664 267338 7676
rect 307386 7664 307392 7676
rect 267332 7636 307392 7664
rect 267332 7624 267338 7636
rect 307386 7624 307392 7636
rect 307444 7624 307450 7676
rect 308858 7624 308864 7676
rect 308916 7664 308922 7676
rect 506014 7664 506020 7676
rect 308916 7636 506020 7664
rect 308916 7624 308922 7636
rect 506014 7624 506020 7636
rect 506072 7624 506078 7676
rect 153930 7556 153936 7608
rect 153988 7596 153994 7608
rect 234982 7596 234988 7608
rect 153988 7568 234988 7596
rect 153988 7556 153994 7568
rect 234982 7556 234988 7568
rect 235040 7556 235046 7608
rect 268746 7556 268752 7608
rect 268804 7596 268810 7608
rect 310974 7596 310980 7608
rect 268804 7568 310980 7596
rect 268804 7556 268810 7568
rect 310974 7556 310980 7568
rect 311032 7556 311038 7608
rect 311618 7556 311624 7608
rect 311676 7596 311682 7608
rect 520366 7596 520372 7608
rect 311676 7568 520372 7596
rect 311676 7556 311682 7568
rect 520366 7556 520372 7568
rect 520424 7556 520430 7608
rect 200390 7488 200396 7540
rect 200448 7528 200454 7540
rect 244826 7528 244832 7540
rect 200448 7500 244832 7528
rect 200448 7488 200454 7500
rect 244826 7488 244832 7500
rect 244884 7488 244890 7540
rect 300762 7488 300768 7540
rect 300820 7528 300826 7540
rect 469122 7528 469128 7540
rect 300820 7500 469128 7528
rect 300820 7488 300826 7500
rect 469122 7488 469128 7500
rect 469180 7488 469186 7540
rect 203886 7420 203892 7472
rect 203944 7460 203950 7472
rect 246022 7460 246028 7472
rect 203944 7432 246028 7460
rect 203944 7420 203950 7432
rect 246022 7420 246028 7432
rect 246080 7420 246086 7472
rect 300670 7420 300676 7472
rect 300728 7460 300734 7472
rect 465626 7460 465632 7472
rect 300728 7432 465632 7460
rect 300728 7420 300734 7432
rect 465626 7420 465632 7432
rect 465684 7420 465690 7472
rect 207474 7352 207480 7404
rect 207532 7392 207538 7404
rect 246390 7392 246396 7404
rect 207532 7364 246396 7392
rect 207532 7352 207538 7364
rect 246390 7352 246396 7364
rect 246448 7352 246454 7404
rect 299382 7352 299388 7404
rect 299440 7392 299446 7404
rect 462038 7392 462044 7404
rect 299440 7364 462044 7392
rect 299440 7352 299446 7364
rect 462038 7352 462044 7364
rect 462096 7352 462102 7404
rect 211062 7284 211068 7336
rect 211120 7324 211126 7336
rect 247402 7324 247408 7336
rect 211120 7296 247408 7324
rect 211120 7284 211126 7296
rect 247402 7284 247408 7296
rect 247460 7284 247466 7336
rect 299290 7284 299296 7336
rect 299348 7324 299354 7336
rect 458450 7324 458456 7336
rect 299348 7296 458456 7324
rect 299348 7284 299354 7296
rect 458450 7284 458456 7296
rect 458508 7284 458514 7336
rect 214650 7216 214656 7268
rect 214708 7256 214714 7268
rect 247494 7256 247500 7268
rect 214708 7228 247500 7256
rect 214708 7216 214714 7228
rect 247494 7216 247500 7228
rect 247552 7216 247558 7268
rect 297910 7216 297916 7268
rect 297968 7256 297974 7268
rect 454862 7256 454868 7268
rect 297968 7228 454868 7256
rect 297968 7216 297974 7228
rect 454862 7216 454868 7228
rect 454920 7216 454926 7268
rect 218146 7148 218152 7200
rect 218204 7188 218210 7200
rect 248782 7188 248788 7200
rect 218204 7160 248788 7188
rect 218204 7148 218210 7160
rect 248782 7148 248788 7160
rect 248840 7148 248846 7200
rect 298002 7148 298008 7200
rect 298060 7188 298066 7200
rect 451366 7188 451372 7200
rect 298060 7160 451372 7188
rect 298060 7148 298066 7160
rect 451366 7148 451372 7160
rect 451424 7148 451430 7200
rect 221734 7080 221740 7132
rect 221792 7120 221798 7132
rect 248690 7120 248696 7132
rect 221792 7092 248696 7120
rect 221792 7080 221798 7092
rect 248690 7080 248696 7092
rect 248748 7080 248754 7132
rect 296530 7080 296536 7132
rect 296588 7120 296594 7132
rect 447778 7120 447784 7132
rect 296588 7092 447784 7120
rect 296588 7080 296594 7092
rect 447778 7080 447784 7092
rect 447836 7080 447842 7132
rect 225322 7012 225328 7064
rect 225380 7052 225386 7064
rect 250254 7052 250260 7064
rect 225380 7024 250260 7052
rect 225380 7012 225386 7024
rect 250254 7012 250260 7024
rect 250312 7012 250318 7064
rect 296622 7012 296628 7064
rect 296680 7052 296686 7064
rect 444190 7052 444196 7064
rect 296680 7024 444196 7052
rect 296680 7012 296686 7024
rect 444190 7012 444196 7024
rect 444248 7012 444254 7064
rect 228910 6944 228916 6996
rect 228968 6984 228974 6996
rect 250162 6984 250168 6996
rect 228968 6956 250168 6984
rect 228968 6944 228974 6956
rect 250162 6944 250168 6956
rect 250220 6944 250226 6996
rect 270126 6944 270132 6996
rect 270184 6984 270190 6996
rect 320450 6984 320456 6996
rect 270184 6956 320456 6984
rect 270184 6944 270190 6956
rect 320450 6944 320456 6956
rect 320508 6944 320514 6996
rect 322474 6944 322480 6996
rect 322532 6984 322538 6996
rect 328454 6984 328460 6996
rect 322532 6956 328460 6984
rect 322532 6944 322538 6956
rect 328454 6944 328460 6956
rect 328512 6944 328518 6996
rect 331490 6944 331496 6996
rect 331548 6984 331554 6996
rect 332410 6984 332416 6996
rect 331548 6956 332416 6984
rect 331548 6944 331554 6956
rect 332410 6944 332416 6956
rect 332468 6944 332474 6996
rect 339678 6944 339684 6996
rect 339736 6984 339742 6996
rect 340690 6984 340696 6996
rect 339736 6956 340696 6984
rect 339736 6944 339742 6956
rect 340690 6944 340696 6956
rect 340748 6944 340754 6996
rect 329098 6876 329104 6928
rect 329156 6916 329162 6928
rect 329190 6916 329196 6928
rect 329156 6888 329196 6916
rect 329156 6876 329162 6888
rect 329190 6876 329196 6888
rect 329248 6876 329254 6928
rect 332962 6876 332968 6928
rect 333020 6916 333026 6928
rect 333146 6916 333152 6928
rect 333020 6888 333152 6916
rect 333020 6876 333026 6888
rect 333146 6876 333152 6888
rect 333204 6876 333210 6928
rect 195606 6808 195612 6860
rect 195664 6848 195670 6860
rect 243078 6848 243084 6860
rect 195664 6820 243084 6848
rect 195664 6808 195670 6820
rect 243078 6808 243084 6820
rect 243136 6808 243142 6860
rect 281350 6808 281356 6860
rect 281408 6848 281414 6860
rect 376386 6848 376392 6860
rect 281408 6820 376392 6848
rect 281408 6808 281414 6820
rect 376386 6808 376392 6820
rect 376444 6808 376450 6860
rect 192018 6740 192024 6792
rect 192076 6780 192082 6792
rect 243446 6780 243452 6792
rect 192076 6752 243452 6780
rect 192076 6740 192082 6752
rect 243446 6740 243452 6752
rect 243504 6740 243510 6792
rect 260558 6740 260564 6792
rect 260616 6780 260622 6792
rect 271690 6780 271696 6792
rect 260616 6752 271696 6780
rect 260616 6740 260622 6752
rect 271690 6740 271696 6752
rect 271748 6740 271754 6792
rect 282822 6740 282828 6792
rect 282880 6780 282886 6792
rect 379974 6780 379980 6792
rect 282880 6752 379980 6780
rect 282880 6740 282886 6752
rect 379974 6740 379980 6752
rect 380032 6740 380038 6792
rect 188430 6672 188436 6724
rect 188488 6712 188494 6724
rect 242158 6712 242164 6724
rect 188488 6684 242164 6712
rect 188488 6672 188494 6684
rect 242158 6672 242164 6684
rect 242216 6672 242222 6724
rect 258810 6672 258816 6724
rect 258868 6712 258874 6724
rect 269298 6712 269304 6724
rect 258868 6684 269304 6712
rect 258868 6672 258874 6684
rect 269298 6672 269304 6684
rect 269356 6672 269362 6724
rect 282730 6672 282736 6724
rect 282788 6712 282794 6724
rect 383562 6712 383568 6724
rect 282788 6684 383568 6712
rect 282788 6672 282794 6684
rect 383562 6672 383568 6684
rect 383620 6672 383626 6724
rect 184842 6604 184848 6656
rect 184900 6644 184906 6656
rect 241790 6644 241796 6656
rect 184900 6616 241796 6644
rect 184900 6604 184906 6616
rect 241790 6604 241796 6616
rect 241848 6604 241854 6656
rect 260466 6604 260472 6656
rect 260524 6644 260530 6656
rect 272886 6644 272892 6656
rect 260524 6616 272892 6644
rect 260524 6604 260530 6616
rect 272886 6604 272892 6616
rect 272944 6604 272950 6656
rect 284202 6604 284208 6656
rect 284260 6644 284266 6656
rect 387058 6644 387064 6656
rect 284260 6616 387064 6644
rect 284260 6604 284266 6616
rect 387058 6604 387064 6616
rect 387116 6604 387122 6656
rect 181346 6536 181352 6588
rect 181404 6576 181410 6588
rect 240410 6576 240416 6588
rect 181404 6548 240416 6576
rect 181404 6536 181410 6548
rect 240410 6536 240416 6548
rect 240468 6536 240474 6588
rect 261846 6536 261852 6588
rect 261904 6576 261910 6588
rect 276474 6576 276480 6588
rect 261904 6548 276480 6576
rect 261904 6536 261910 6548
rect 276474 6536 276480 6548
rect 276532 6536 276538 6588
rect 285490 6536 285496 6588
rect 285548 6576 285554 6588
rect 390646 6576 390652 6588
rect 285548 6548 390652 6576
rect 285548 6536 285554 6548
rect 390646 6536 390652 6548
rect 390704 6536 390710 6588
rect 177758 6468 177764 6520
rect 177816 6508 177822 6520
rect 240318 6508 240324 6520
rect 177816 6480 240324 6508
rect 177816 6468 177822 6480
rect 240318 6468 240324 6480
rect 240376 6468 240382 6520
rect 260374 6468 260380 6520
rect 260432 6508 260438 6520
rect 275278 6508 275284 6520
rect 260432 6480 275284 6508
rect 260432 6468 260438 6480
rect 275278 6468 275284 6480
rect 275336 6468 275342 6520
rect 285582 6468 285588 6520
rect 285640 6508 285646 6520
rect 394234 6508 394240 6520
rect 285640 6480 394240 6508
rect 285640 6468 285646 6480
rect 394234 6468 394240 6480
rect 394292 6468 394298 6520
rect 174170 6400 174176 6452
rect 174228 6440 174234 6452
rect 238846 6440 238852 6452
rect 174228 6412 238852 6440
rect 174228 6400 174234 6412
rect 238846 6400 238852 6412
rect 238904 6400 238910 6452
rect 261754 6400 261760 6452
rect 261812 6440 261818 6452
rect 278866 6440 278872 6452
rect 261812 6412 278872 6440
rect 261812 6400 261818 6412
rect 278866 6400 278872 6412
rect 278924 6400 278930 6452
rect 286870 6400 286876 6452
rect 286928 6440 286934 6452
rect 397822 6440 397828 6452
rect 286928 6412 397828 6440
rect 286928 6400 286934 6412
rect 397822 6400 397828 6412
rect 397880 6400 397886 6452
rect 170582 6332 170588 6384
rect 170640 6372 170646 6384
rect 238938 6372 238944 6384
rect 170640 6344 238944 6372
rect 170640 6332 170646 6344
rect 238938 6332 238944 6344
rect 238996 6332 239002 6384
rect 261662 6332 261668 6384
rect 261720 6372 261726 6384
rect 280065 6375 280123 6381
rect 280065 6372 280077 6375
rect 261720 6344 280077 6372
rect 261720 6332 261726 6344
rect 280065 6341 280077 6344
rect 280111 6341 280123 6375
rect 280065 6335 280123 6341
rect 286962 6332 286968 6384
rect 287020 6372 287026 6384
rect 401318 6372 401324 6384
rect 287020 6344 401324 6372
rect 287020 6332 287026 6344
rect 401318 6332 401324 6344
rect 401376 6332 401382 6384
rect 159910 6264 159916 6316
rect 159968 6304 159974 6316
rect 236178 6304 236184 6316
rect 159968 6276 236184 6304
rect 159968 6264 159974 6276
rect 236178 6264 236184 6276
rect 236236 6264 236242 6316
rect 261938 6264 261944 6316
rect 261996 6304 262002 6316
rect 282454 6304 282460 6316
rect 261996 6276 282460 6304
rect 261996 6264 262002 6276
rect 282454 6264 282460 6276
rect 282512 6264 282518 6316
rect 288342 6264 288348 6316
rect 288400 6304 288406 6316
rect 404906 6304 404912 6316
rect 288400 6276 404912 6304
rect 288400 6264 288406 6276
rect 404906 6264 404912 6276
rect 404964 6264 404970 6316
rect 156322 6196 156328 6248
rect 156380 6236 156386 6248
rect 236086 6236 236092 6248
rect 156380 6208 236092 6236
rect 156380 6196 156386 6208
rect 236086 6196 236092 6208
rect 236144 6196 236150 6248
rect 262950 6196 262956 6248
rect 263008 6236 263014 6248
rect 285950 6236 285956 6248
rect 263008 6208 285956 6236
rect 263008 6196 263014 6208
rect 285950 6196 285956 6208
rect 286008 6196 286014 6248
rect 288250 6196 288256 6248
rect 288308 6236 288314 6248
rect 408586 6236 408592 6248
rect 288308 6208 408592 6236
rect 288308 6196 288314 6208
rect 408586 6196 408592 6208
rect 408644 6196 408650 6248
rect 152734 6128 152740 6180
rect 152792 6168 152798 6180
rect 235258 6168 235264 6180
rect 152792 6140 235264 6168
rect 152792 6128 152798 6140
rect 235258 6128 235264 6140
rect 235316 6128 235322 6180
rect 263134 6128 263140 6180
rect 263192 6168 263198 6180
rect 289538 6168 289544 6180
rect 263192 6140 289544 6168
rect 263192 6128 263198 6140
rect 289538 6128 289544 6140
rect 289596 6128 289602 6180
rect 289722 6128 289728 6180
rect 289780 6168 289786 6180
rect 412082 6168 412088 6180
rect 289780 6140 412088 6168
rect 289780 6128 289786 6140
rect 412082 6128 412088 6140
rect 412140 6128 412146 6180
rect 199194 6060 199200 6112
rect 199252 6100 199258 6112
rect 244734 6100 244740 6112
rect 199252 6072 244740 6100
rect 199252 6060 199258 6072
rect 244734 6060 244740 6072
rect 244792 6060 244798 6112
rect 281442 6060 281448 6112
rect 281500 6100 281506 6112
rect 372798 6100 372804 6112
rect 281500 6072 372804 6100
rect 281500 6060 281506 6072
rect 372798 6060 372804 6072
rect 372856 6060 372862 6112
rect 202690 5992 202696 6044
rect 202748 6032 202754 6044
rect 245654 6032 245660 6044
rect 202748 6004 245660 6032
rect 202748 5992 202754 6004
rect 245654 5992 245660 6004
rect 245712 5992 245718 6044
rect 279970 5992 279976 6044
rect 280028 6032 280034 6044
rect 369210 6032 369216 6044
rect 280028 6004 369216 6032
rect 280028 5992 280034 6004
rect 369210 5992 369216 6004
rect 369268 5992 369274 6044
rect 206278 5924 206284 5976
rect 206336 5964 206342 5976
rect 245930 5964 245936 5976
rect 206336 5936 245936 5964
rect 206336 5924 206342 5936
rect 245930 5924 245936 5936
rect 245988 5924 245994 5976
rect 280062 5924 280068 5976
rect 280120 5964 280126 5976
rect 365714 5964 365720 5976
rect 280120 5936 365720 5964
rect 280120 5924 280126 5936
rect 365714 5924 365720 5936
rect 365772 5924 365778 5976
rect 209866 5856 209872 5908
rect 209924 5896 209930 5908
rect 247218 5896 247224 5908
rect 209924 5868 247224 5896
rect 209924 5856 209930 5868
rect 247218 5856 247224 5868
rect 247276 5856 247282 5908
rect 278682 5856 278688 5908
rect 278740 5896 278746 5908
rect 362126 5896 362132 5908
rect 278740 5868 362132 5896
rect 278740 5856 278746 5868
rect 362126 5856 362132 5868
rect 362184 5856 362190 5908
rect 213454 5788 213460 5840
rect 213512 5828 213518 5840
rect 247678 5828 247684 5840
rect 213512 5800 247684 5828
rect 213512 5788 213518 5800
rect 247678 5788 247684 5800
rect 247736 5788 247742 5840
rect 278590 5788 278596 5840
rect 278648 5828 278654 5840
rect 358538 5828 358544 5840
rect 278648 5800 358544 5828
rect 278648 5788 278654 5800
rect 358538 5788 358544 5800
rect 358596 5788 358602 5840
rect 217042 5720 217048 5772
rect 217100 5760 217106 5772
rect 248598 5760 248604 5772
rect 217100 5732 248604 5760
rect 217100 5720 217106 5732
rect 248598 5720 248604 5732
rect 248656 5720 248662 5772
rect 277210 5720 277216 5772
rect 277268 5760 277274 5772
rect 354950 5760 354956 5772
rect 277268 5732 354956 5760
rect 277268 5720 277274 5732
rect 354950 5720 354956 5732
rect 355008 5720 355014 5772
rect 220538 5652 220544 5704
rect 220596 5692 220602 5704
rect 248506 5692 248512 5704
rect 220596 5664 248512 5692
rect 220596 5652 220602 5664
rect 248506 5652 248512 5664
rect 248564 5652 248570 5704
rect 277302 5652 277308 5704
rect 277360 5692 277366 5704
rect 351362 5692 351368 5704
rect 277360 5664 351368 5692
rect 277360 5652 277366 5664
rect 351362 5652 351368 5664
rect 351420 5652 351426 5704
rect 224126 5584 224132 5636
rect 224184 5624 224190 5636
rect 250070 5624 250076 5636
rect 224184 5596 250076 5624
rect 224184 5584 224190 5596
rect 250070 5584 250076 5596
rect 250128 5584 250134 5636
rect 275554 5584 275560 5636
rect 275612 5624 275618 5636
rect 347866 5624 347872 5636
rect 275612 5596 347872 5624
rect 275612 5584 275618 5596
rect 347866 5584 347872 5596
rect 347924 5584 347930 5636
rect 227714 5516 227720 5568
rect 227772 5556 227778 5568
rect 249978 5556 249984 5568
rect 227772 5528 249984 5556
rect 227772 5516 227778 5528
rect 249978 5516 249984 5528
rect 250036 5516 250042 5568
rect 250257 5559 250315 5565
rect 250257 5525 250269 5559
rect 250303 5556 250315 5559
rect 252646 5556 252652 5568
rect 250303 5528 252652 5556
rect 250303 5525 250315 5528
rect 250257 5519 250315 5525
rect 252646 5516 252652 5528
rect 252704 5516 252710 5568
rect 267277 5559 267335 5565
rect 267277 5525 267289 5559
rect 267323 5556 267335 5559
rect 268381 5559 268439 5565
rect 268381 5556 268393 5559
rect 267323 5528 268393 5556
rect 267323 5525 267335 5528
rect 267277 5519 267335 5525
rect 268381 5525 268393 5528
rect 268427 5525 268439 5559
rect 268381 5519 268439 5525
rect 275922 5516 275928 5568
rect 275980 5556 275986 5568
rect 344278 5556 344284 5568
rect 275980 5528 344284 5556
rect 275980 5516 275986 5528
rect 344278 5516 344284 5528
rect 344336 5516 344342 5568
rect 124214 5448 124220 5500
rect 124272 5488 124278 5500
rect 191098 5488 191104 5500
rect 124272 5460 191104 5488
rect 124272 5448 124278 5460
rect 191098 5448 191104 5460
rect 191156 5448 191162 5500
rect 194410 5448 194416 5500
rect 194468 5488 194474 5500
rect 243078 5488 243084 5500
rect 194468 5460 243084 5488
rect 194468 5448 194474 5460
rect 243078 5448 243084 5460
rect 243136 5448 243142 5500
rect 243170 5448 243176 5500
rect 243228 5488 243234 5500
rect 254026 5488 254032 5500
rect 243228 5460 254032 5488
rect 243228 5448 243234 5460
rect 254026 5448 254032 5460
rect 254084 5448 254090 5500
rect 255038 5448 255044 5500
rect 255096 5488 255102 5500
rect 255774 5488 255780 5500
rect 255096 5460 255780 5488
rect 255096 5448 255102 5460
rect 255774 5448 255780 5460
rect 255832 5448 255838 5500
rect 256234 5448 256240 5500
rect 256292 5488 256298 5500
rect 257246 5488 257252 5500
rect 256292 5460 257252 5488
rect 256292 5448 256298 5460
rect 257246 5448 257252 5460
rect 257304 5448 257310 5500
rect 257798 5448 257804 5500
rect 257856 5488 257862 5500
rect 258626 5488 258632 5500
rect 257856 5460 258632 5488
rect 257856 5448 257862 5460
rect 258626 5448 258632 5460
rect 258684 5448 258690 5500
rect 264882 5448 264888 5500
rect 264940 5488 264946 5500
rect 291930 5488 291936 5500
rect 264940 5460 291936 5488
rect 264940 5448 264946 5460
rect 291930 5448 291936 5460
rect 291988 5448 291994 5500
rect 311710 5448 311716 5500
rect 311768 5488 311774 5500
rect 522666 5488 522672 5500
rect 311768 5460 522672 5488
rect 311768 5448 311774 5460
rect 522666 5448 522672 5460
rect 522724 5448 522730 5500
rect 113542 5380 113548 5432
rect 113600 5420 113606 5432
rect 182818 5420 182824 5432
rect 113600 5392 182824 5420
rect 113600 5380 113606 5392
rect 182818 5380 182824 5392
rect 182876 5380 182882 5432
rect 187234 5380 187240 5432
rect 187292 5420 187298 5432
rect 241606 5420 241612 5432
rect 187292 5392 241612 5420
rect 187292 5380 187298 5392
rect 241606 5380 241612 5392
rect 241664 5380 241670 5432
rect 241974 5380 241980 5432
rect 242032 5420 242038 5432
rect 252925 5423 252983 5429
rect 252925 5420 252937 5423
rect 242032 5392 252937 5420
rect 242032 5380 242038 5392
rect 252925 5389 252937 5392
rect 252971 5389 252983 5423
rect 252925 5383 252983 5389
rect 257706 5380 257712 5432
rect 257764 5420 257770 5432
rect 259822 5420 259828 5432
rect 257764 5392 259828 5420
rect 257764 5380 257770 5392
rect 259822 5380 259828 5392
rect 259880 5380 259886 5432
rect 264698 5380 264704 5432
rect 264756 5420 264762 5432
rect 294322 5420 294328 5432
rect 264756 5392 294328 5420
rect 264756 5380 264762 5392
rect 294322 5380 294328 5392
rect 294380 5380 294386 5432
rect 313090 5380 313096 5432
rect 313148 5420 313154 5432
rect 526254 5420 526260 5432
rect 313148 5392 526260 5420
rect 313148 5380 313154 5392
rect 526254 5380 526260 5392
rect 526312 5380 526318 5432
rect 125410 5312 125416 5364
rect 125468 5352 125474 5364
rect 195238 5352 195244 5364
rect 125468 5324 195244 5352
rect 125468 5312 125474 5324
rect 195238 5312 195244 5324
rect 195296 5312 195302 5364
rect 197998 5312 198004 5364
rect 198056 5352 198062 5364
rect 244366 5352 244372 5364
rect 198056 5324 244372 5352
rect 198056 5312 198062 5324
rect 244366 5312 244372 5324
rect 244424 5312 244430 5364
rect 244642 5312 244648 5364
rect 244700 5352 244706 5364
rect 254394 5352 254400 5364
rect 244700 5324 254400 5352
rect 244700 5312 244706 5324
rect 254394 5312 254400 5324
rect 254452 5312 254458 5364
rect 257982 5312 257988 5364
rect 258040 5352 258046 5364
rect 261018 5352 261024 5364
rect 258040 5324 261024 5352
rect 258040 5312 258046 5324
rect 261018 5312 261024 5324
rect 261076 5312 261082 5364
rect 264606 5312 264612 5364
rect 264664 5352 264670 5364
rect 267277 5355 267335 5361
rect 267277 5352 267289 5355
rect 264664 5324 267289 5352
rect 264664 5312 264670 5324
rect 267277 5321 267289 5324
rect 267323 5321 267335 5355
rect 267277 5315 267335 5321
rect 267366 5312 267372 5364
rect 267424 5352 267430 5364
rect 268289 5355 268347 5361
rect 268289 5352 268301 5355
rect 267424 5324 268301 5352
rect 267424 5312 267430 5324
rect 268289 5321 268301 5324
rect 268335 5321 268347 5355
rect 268289 5315 268347 5321
rect 268381 5355 268439 5361
rect 268381 5321 268393 5355
rect 268427 5352 268439 5355
rect 295518 5352 295524 5364
rect 268427 5324 295524 5352
rect 268427 5321 268439 5324
rect 268381 5315 268439 5321
rect 295518 5312 295524 5324
rect 295576 5312 295582 5364
rect 313182 5312 313188 5364
rect 313240 5352 313246 5364
rect 529842 5352 529848 5364
rect 313240 5324 529848 5352
rect 313240 5312 313246 5324
rect 529842 5312 529848 5324
rect 529900 5312 529906 5364
rect 158714 5244 158720 5296
rect 158772 5284 158778 5296
rect 235902 5284 235908 5296
rect 158772 5256 235908 5284
rect 158772 5244 158778 5256
rect 235902 5244 235908 5256
rect 235960 5244 235966 5296
rect 235994 5244 236000 5296
rect 236052 5284 236058 5296
rect 251450 5284 251456 5296
rect 236052 5256 251456 5284
rect 236052 5244 236058 5256
rect 251450 5244 251456 5256
rect 251508 5244 251514 5296
rect 257890 5244 257896 5296
rect 257948 5284 257954 5296
rect 262214 5284 262220 5296
rect 257948 5256 262220 5284
rect 257948 5244 257954 5256
rect 262214 5244 262220 5256
rect 262272 5244 262278 5296
rect 266078 5244 266084 5296
rect 266136 5284 266142 5296
rect 297910 5284 297916 5296
rect 266136 5256 297916 5284
rect 266136 5244 266142 5256
rect 297910 5244 297916 5256
rect 297968 5244 297974 5296
rect 314470 5244 314476 5296
rect 314528 5284 314534 5296
rect 533430 5284 533436 5296
rect 314528 5256 533436 5284
rect 314528 5244 314534 5256
rect 533430 5244 533436 5256
rect 533488 5244 533494 5296
rect 155126 5176 155132 5228
rect 155184 5216 155190 5228
rect 235166 5216 235172 5228
rect 155184 5188 235172 5216
rect 155184 5176 155190 5188
rect 235166 5176 235172 5188
rect 235224 5176 235230 5228
rect 238386 5176 238392 5228
rect 238444 5216 238450 5228
rect 252830 5216 252836 5228
rect 238444 5188 252836 5216
rect 238444 5176 238450 5188
rect 252830 5176 252836 5188
rect 252888 5176 252894 5228
rect 266170 5176 266176 5228
rect 266228 5216 266234 5228
rect 299106 5216 299112 5228
rect 266228 5188 299112 5216
rect 266228 5176 266234 5188
rect 299106 5176 299112 5188
rect 299164 5176 299170 5228
rect 314378 5176 314384 5228
rect 314436 5216 314442 5228
rect 536926 5216 536932 5228
rect 314436 5188 536932 5216
rect 314436 5176 314442 5188
rect 536926 5176 536932 5188
rect 536984 5176 536990 5228
rect 151538 5108 151544 5160
rect 151596 5148 151602 5160
rect 234706 5148 234712 5160
rect 151596 5120 234712 5148
rect 151596 5108 151602 5120
rect 234706 5108 234712 5120
rect 234764 5108 234770 5160
rect 237190 5108 237196 5160
rect 237248 5148 237254 5160
rect 252738 5148 252744 5160
rect 237248 5120 252744 5148
rect 237248 5108 237254 5120
rect 252738 5108 252744 5120
rect 252796 5108 252802 5160
rect 266262 5108 266268 5160
rect 266320 5148 266326 5160
rect 301406 5148 301412 5160
rect 266320 5120 301412 5148
rect 266320 5108 266326 5120
rect 301406 5108 301412 5120
rect 301464 5108 301470 5160
rect 315850 5108 315856 5160
rect 315908 5148 315914 5160
rect 540514 5148 540520 5160
rect 315908 5120 540520 5148
rect 315908 5108 315914 5120
rect 540514 5108 540520 5120
rect 540572 5108 540578 5160
rect 148042 5040 148048 5092
rect 148100 5080 148106 5092
rect 233326 5080 233332 5092
rect 148100 5052 233332 5080
rect 148100 5040 148106 5052
rect 233326 5040 233332 5052
rect 233384 5040 233390 5092
rect 234798 5040 234804 5092
rect 234856 5080 234862 5092
rect 251634 5080 251640 5092
rect 234856 5052 251640 5080
rect 234856 5040 234862 5052
rect 251634 5040 251640 5052
rect 251692 5040 251698 5092
rect 267642 5040 267648 5092
rect 267700 5080 267706 5092
rect 270681 5083 270739 5089
rect 267700 5052 270632 5080
rect 267700 5040 267706 5052
rect 144454 4972 144460 5024
rect 144512 5012 144518 5024
rect 233234 5012 233240 5024
rect 144512 4984 233240 5012
rect 144512 4972 144518 4984
rect 233234 4972 233240 4984
rect 233292 4972 233298 5024
rect 233694 4972 233700 5024
rect 233752 5012 233758 5024
rect 251358 5012 251364 5024
rect 233752 4984 251364 5012
rect 233752 4972 233758 4984
rect 251358 4972 251364 4984
rect 251416 4972 251422 5024
rect 260742 4972 260748 5024
rect 260800 5012 260806 5024
rect 270494 5012 270500 5024
rect 260800 4984 270500 5012
rect 260800 4972 260806 4984
rect 270494 4972 270500 4984
rect 270552 4972 270558 5024
rect 270604 5012 270632 5052
rect 270681 5049 270693 5083
rect 270727 5080 270739 5083
rect 302602 5080 302608 5092
rect 270727 5052 302608 5080
rect 270727 5049 270739 5052
rect 270681 5043 270739 5049
rect 302602 5040 302608 5052
rect 302660 5040 302666 5092
rect 315942 5040 315948 5092
rect 316000 5080 316006 5092
rect 544102 5080 544108 5092
rect 316000 5052 544108 5080
rect 316000 5040 316006 5052
rect 544102 5040 544108 5052
rect 544160 5040 544166 5092
rect 304994 5012 305000 5024
rect 270604 4984 305000 5012
rect 304994 4972 305000 4984
rect 305052 4972 305058 5024
rect 317322 4972 317328 5024
rect 317380 5012 317386 5024
rect 547690 5012 547696 5024
rect 317380 4984 547696 5012
rect 317380 4972 317386 4984
rect 547690 4972 547696 4984
rect 547748 4972 547754 5024
rect 140866 4904 140872 4956
rect 140924 4944 140930 4956
rect 232406 4944 232412 4956
rect 140924 4916 232412 4944
rect 140924 4904 140930 4916
rect 232406 4904 232412 4916
rect 232464 4904 232470 4956
rect 232498 4904 232504 4956
rect 232556 4944 232562 4956
rect 251726 4944 251732 4956
rect 232556 4916 251732 4944
rect 232556 4904 232562 4916
rect 251726 4904 251732 4916
rect 251784 4904 251790 4956
rect 259270 4904 259276 4956
rect 259328 4944 259334 4956
rect 268102 4944 268108 4956
rect 259328 4916 268108 4944
rect 259328 4904 259334 4916
rect 268102 4904 268108 4916
rect 268160 4904 268166 4956
rect 268289 4947 268347 4953
rect 268289 4913 268301 4947
rect 268335 4944 268347 4947
rect 306190 4944 306196 4956
rect 268335 4916 306196 4944
rect 268335 4913 268347 4916
rect 268289 4907 268347 4913
rect 306190 4904 306196 4916
rect 306248 4904 306254 4956
rect 318610 4904 318616 4956
rect 318668 4944 318674 4956
rect 551186 4944 551192 4956
rect 318668 4916 551192 4944
rect 318668 4904 318674 4916
rect 551186 4904 551192 4916
rect 551244 4904 551250 4956
rect 133782 4836 133788 4888
rect 133840 4876 133846 4888
rect 231026 4876 231032 4888
rect 133840 4848 231032 4876
rect 133840 4836 133846 4848
rect 231026 4836 231032 4848
rect 231084 4836 231090 4888
rect 231302 4836 231308 4888
rect 231360 4876 231366 4888
rect 251542 4876 251548 4888
rect 231360 4848 251548 4876
rect 231360 4836 231366 4848
rect 251542 4836 251548 4848
rect 251600 4836 251606 4888
rect 262122 4836 262128 4888
rect 262180 4876 262186 4888
rect 267369 4879 267427 4885
rect 267369 4876 267381 4879
rect 262180 4848 267381 4876
rect 262180 4836 262186 4848
rect 267369 4845 267381 4848
rect 267415 4845 267427 4879
rect 267369 4839 267427 4845
rect 267458 4836 267464 4888
rect 267516 4876 267522 4888
rect 308582 4876 308588 4888
rect 267516 4848 308588 4876
rect 267516 4836 267522 4848
rect 308582 4836 308588 4848
rect 308640 4836 308646 4888
rect 318702 4836 318708 4888
rect 318760 4876 318766 4888
rect 554774 4876 554780 4888
rect 318760 4848 554780 4876
rect 318760 4836 318766 4848
rect 554774 4836 554780 4848
rect 554832 4836 554838 4888
rect 127802 4768 127808 4820
rect 127860 4808 127866 4820
rect 229186 4808 229192 4820
rect 127860 4780 229192 4808
rect 127860 4768 127866 4780
rect 229186 4768 229192 4780
rect 229244 4768 229250 4820
rect 230106 4768 230112 4820
rect 230164 4808 230170 4820
rect 251174 4808 251180 4820
rect 230164 4780 251180 4808
rect 230164 4768 230170 4780
rect 251174 4768 251180 4780
rect 251232 4768 251238 4820
rect 262030 4768 262036 4820
rect 262088 4808 262094 4820
rect 264977 4811 265035 4817
rect 264977 4808 264989 4811
rect 262088 4780 264989 4808
rect 262088 4768 262094 4780
rect 264977 4777 264989 4780
rect 265023 4777 265035 4811
rect 264977 4771 265035 4777
rect 265986 4768 265992 4820
rect 266044 4808 266050 4820
rect 266044 4780 268516 4808
rect 266044 4768 266050 4780
rect 106366 4700 106372 4752
rect 106424 4740 106430 4752
rect 106424 4712 118648 4740
rect 106424 4700 106430 4712
rect 118620 4672 118648 4712
rect 120626 4700 120632 4752
rect 120684 4740 120690 4752
rect 135257 4743 135315 4749
rect 135257 4740 135269 4743
rect 120684 4712 135269 4740
rect 120684 4700 120690 4712
rect 135257 4709 135269 4712
rect 135303 4709 135315 4743
rect 135257 4703 135315 4709
rect 135441 4743 135499 4749
rect 135441 4709 135453 4743
rect 135487 4740 135499 4743
rect 154577 4743 154635 4749
rect 154577 4740 154589 4743
rect 135487 4712 154589 4740
rect 135487 4709 135499 4712
rect 135441 4703 135499 4709
rect 154577 4709 154589 4712
rect 154623 4709 154635 4743
rect 154577 4703 154635 4709
rect 154761 4743 154819 4749
rect 154761 4709 154773 4743
rect 154807 4740 154819 4743
rect 186958 4740 186964 4752
rect 154807 4712 186964 4740
rect 154807 4709 154819 4712
rect 154761 4703 154819 4709
rect 186958 4700 186964 4712
rect 187016 4700 187022 4752
rect 201494 4700 201500 4752
rect 201552 4740 201558 4752
rect 244274 4740 244280 4752
rect 201552 4712 244280 4740
rect 201552 4700 201558 4712
rect 244274 4700 244280 4712
rect 244332 4700 244338 4752
rect 245562 4700 245568 4752
rect 245620 4740 245626 4752
rect 254302 4740 254308 4752
rect 245620 4712 254308 4740
rect 245620 4700 245626 4712
rect 254302 4700 254308 4712
rect 254360 4700 254366 4752
rect 260650 4700 260656 4752
rect 260708 4740 260714 4752
rect 268381 4743 268439 4749
rect 268381 4740 268393 4743
rect 260708 4712 268393 4740
rect 260708 4700 260714 4712
rect 268381 4709 268393 4712
rect 268427 4709 268439 4743
rect 268488 4740 268516 4780
rect 268930 4768 268936 4820
rect 268988 4808 268994 4820
rect 312170 4808 312176 4820
rect 268988 4780 312176 4808
rect 268988 4768 268994 4780
rect 312170 4768 312176 4780
rect 312228 4768 312234 4820
rect 320082 4768 320088 4820
rect 320140 4808 320146 4820
rect 558362 4808 558368 4820
rect 320140 4780 558368 4808
rect 320140 4768 320146 4780
rect 558362 4768 558368 4780
rect 558420 4768 558426 4820
rect 270681 4743 270739 4749
rect 270681 4740 270693 4743
rect 268488 4712 270693 4740
rect 268381 4703 268439 4709
rect 270681 4709 270693 4712
rect 270727 4709 270739 4743
rect 270681 4703 270739 4709
rect 270773 4743 270831 4749
rect 270773 4709 270785 4743
rect 270819 4740 270831 4743
rect 290734 4740 290740 4752
rect 270819 4712 290740 4740
rect 270819 4709 270831 4712
rect 270773 4703 270831 4709
rect 290734 4700 290740 4712
rect 290792 4700 290798 4752
rect 311802 4700 311808 4752
rect 311860 4740 311866 4752
rect 519078 4740 519084 4752
rect 311860 4712 519084 4740
rect 311860 4700 311866 4712
rect 519078 4700 519084 4712
rect 519136 4700 519142 4752
rect 135165 4675 135223 4681
rect 118620 4644 118924 4672
rect 118896 4604 118924 4644
rect 135165 4641 135177 4675
rect 135211 4672 135223 4675
rect 135349 4675 135407 4681
rect 135349 4672 135361 4675
rect 135211 4644 135361 4672
rect 135211 4641 135223 4644
rect 135165 4635 135223 4641
rect 135349 4641 135361 4644
rect 135395 4641 135407 4675
rect 135349 4635 135407 4641
rect 154485 4675 154543 4681
rect 154485 4641 154497 4675
rect 154531 4672 154543 4675
rect 154531 4644 154620 4672
rect 154531 4641 154543 4644
rect 154485 4635 154543 4641
rect 154592 4613 154620 4644
rect 172974 4632 172980 4684
rect 173032 4672 173038 4684
rect 239398 4672 239404 4684
rect 173032 4644 239404 4672
rect 173032 4632 173038 4644
rect 239398 4632 239404 4644
rect 239456 4632 239462 4684
rect 239582 4632 239588 4684
rect 239640 4672 239646 4684
rect 252554 4672 252560 4684
rect 239640 4644 252560 4672
rect 239640 4632 239646 4644
rect 252554 4632 252560 4644
rect 252612 4632 252618 4684
rect 263410 4632 263416 4684
rect 263468 4672 263474 4684
rect 287146 4672 287152 4684
rect 263468 4644 287152 4672
rect 263468 4632 263474 4644
rect 287146 4632 287152 4644
rect 287204 4632 287210 4684
rect 310330 4632 310336 4684
rect 310388 4672 310394 4684
rect 515582 4672 515588 4684
rect 310388 4644 515588 4672
rect 310388 4632 310394 4644
rect 515582 4632 515588 4644
rect 515640 4632 515646 4684
rect 125597 4607 125655 4613
rect 125597 4604 125609 4607
rect 118896 4576 125609 4604
rect 125597 4573 125609 4576
rect 125643 4573 125655 4607
rect 154577 4607 154635 4613
rect 125597 4567 125655 4573
rect 144840 4576 144960 4604
rect 135349 4539 135407 4545
rect 135349 4505 135361 4539
rect 135395 4536 135407 4539
rect 144840 4536 144868 4576
rect 144932 4545 144960 4576
rect 154577 4573 154589 4607
rect 154623 4573 154635 4607
rect 154577 4567 154635 4573
rect 180150 4564 180156 4616
rect 180208 4604 180214 4616
rect 238757 4607 238815 4613
rect 238757 4604 238769 4607
rect 180208 4576 238769 4604
rect 180208 4564 180214 4576
rect 238757 4573 238769 4576
rect 238803 4573 238815 4607
rect 238757 4567 238815 4573
rect 238846 4564 238852 4616
rect 238904 4604 238910 4616
rect 239677 4607 239735 4613
rect 238904 4576 239536 4604
rect 238904 4564 238910 4576
rect 135395 4508 144868 4536
rect 144917 4539 144975 4545
rect 135395 4505 135407 4508
rect 135349 4499 135407 4505
rect 144917 4505 144929 4539
rect 144963 4505 144975 4539
rect 144917 4499 144975 4505
rect 164145 4539 164203 4545
rect 164145 4505 164157 4539
rect 164191 4536 164203 4539
rect 173158 4536 173164 4548
rect 164191 4508 173164 4536
rect 164191 4505 164203 4508
rect 164145 4499 164203 4505
rect 173158 4496 173164 4508
rect 173216 4496 173222 4548
rect 208670 4496 208676 4548
rect 208728 4536 208734 4548
rect 239033 4539 239091 4545
rect 208728 4508 238984 4536
rect 208728 4496 208734 4508
rect 125597 4471 125655 4477
rect 125597 4437 125609 4471
rect 125643 4468 125655 4471
rect 135165 4471 135223 4477
rect 135165 4468 135177 4471
rect 125643 4440 135177 4468
rect 125643 4437 125655 4440
rect 125597 4431 125655 4437
rect 135165 4437 135177 4440
rect 135211 4437 135223 4471
rect 135165 4431 135223 4437
rect 212258 4428 212264 4480
rect 212316 4468 212322 4480
rect 238846 4468 238852 4480
rect 212316 4440 238852 4468
rect 212316 4428 212322 4440
rect 238846 4428 238852 4440
rect 238904 4428 238910 4480
rect 238956 4468 238984 4508
rect 239033 4505 239045 4539
rect 239079 4536 239091 4539
rect 239401 4539 239459 4545
rect 239401 4536 239413 4539
rect 239079 4508 239413 4536
rect 239079 4505 239091 4508
rect 239033 4499 239091 4505
rect 239401 4505 239413 4508
rect 239447 4505 239459 4539
rect 239508 4536 239536 4576
rect 239677 4573 239689 4607
rect 239723 4604 239735 4607
rect 240594 4604 240600 4616
rect 239723 4576 240600 4604
rect 239723 4573 239735 4576
rect 239677 4567 239735 4573
rect 240594 4564 240600 4576
rect 240652 4564 240658 4616
rect 240778 4564 240784 4616
rect 240836 4604 240842 4616
rect 246669 4607 246727 4613
rect 246669 4604 246681 4607
rect 240836 4576 246681 4604
rect 240836 4564 240842 4576
rect 246669 4573 246681 4576
rect 246715 4573 246727 4607
rect 246669 4567 246727 4573
rect 246758 4564 246764 4616
rect 246816 4604 246822 4616
rect 254578 4604 254584 4616
rect 246816 4576 254584 4604
rect 246816 4564 246822 4576
rect 254578 4564 254584 4576
rect 254636 4564 254642 4616
rect 263318 4564 263324 4616
rect 263376 4604 263382 4616
rect 288342 4604 288348 4616
rect 263376 4576 288348 4604
rect 263376 4564 263382 4576
rect 288342 4564 288348 4576
rect 288400 4564 288406 4616
rect 310422 4564 310428 4616
rect 310480 4604 310486 4616
rect 511994 4604 512000 4616
rect 310480 4576 512000 4604
rect 310480 4564 310486 4576
rect 511994 4564 512000 4576
rect 512052 4564 512058 4616
rect 247586 4536 247592 4548
rect 239508 4508 247592 4536
rect 239401 4499 239459 4505
rect 247586 4496 247592 4508
rect 247644 4496 247650 4548
rect 247954 4496 247960 4548
rect 248012 4536 248018 4548
rect 254118 4536 254124 4548
rect 248012 4508 254124 4536
rect 248012 4496 248018 4508
rect 254118 4496 254124 4508
rect 254176 4496 254182 4548
rect 259086 4496 259092 4548
rect 259144 4536 259150 4548
rect 263413 4539 263471 4545
rect 263413 4536 263425 4539
rect 259144 4508 263425 4536
rect 259144 4496 259150 4508
rect 263413 4505 263425 4508
rect 263459 4505 263471 4539
rect 263413 4499 263471 4505
rect 263502 4496 263508 4548
rect 263560 4536 263566 4548
rect 284754 4536 284760 4548
rect 263560 4508 284760 4536
rect 263560 4496 263566 4508
rect 284754 4496 284760 4508
rect 284812 4496 284818 4548
rect 309042 4496 309048 4548
rect 309100 4536 309106 4548
rect 508406 4536 508412 4548
rect 309100 4508 508412 4536
rect 309100 4496 309106 4508
rect 508406 4496 508412 4508
rect 508464 4496 508470 4548
rect 246206 4468 246212 4480
rect 238956 4440 246212 4468
rect 246206 4428 246212 4440
rect 246264 4428 246270 4480
rect 246669 4471 246727 4477
rect 246669 4437 246681 4471
rect 246715 4468 246727 4471
rect 250257 4471 250315 4477
rect 250257 4468 250269 4471
rect 246715 4440 250269 4468
rect 246715 4437 246727 4440
rect 246669 4431 246727 4437
rect 250257 4437 250269 4440
rect 250303 4437 250315 4471
rect 250257 4431 250315 4437
rect 250346 4428 250352 4480
rect 250404 4468 250410 4480
rect 255314 4468 255320 4480
rect 250404 4440 255320 4468
rect 250404 4428 250410 4440
rect 255314 4428 255320 4440
rect 255372 4428 255378 4480
rect 263226 4428 263232 4480
rect 263284 4468 263290 4480
rect 283650 4468 283656 4480
rect 263284 4440 283656 4468
rect 263284 4428 263290 4440
rect 283650 4428 283656 4440
rect 283708 4428 283714 4480
rect 308950 4428 308956 4480
rect 309008 4468 309014 4480
rect 504818 4468 504824 4480
rect 309008 4440 504824 4468
rect 309008 4428 309014 4440
rect 504818 4428 504824 4440
rect 504876 4428 504882 4480
rect 144917 4403 144975 4409
rect 144917 4369 144929 4403
rect 144963 4400 144975 4403
rect 154485 4403 154543 4409
rect 154485 4400 154497 4403
rect 144963 4372 154497 4400
rect 144963 4369 144975 4372
rect 144917 4363 144975 4369
rect 154485 4369 154497 4372
rect 154531 4369 154543 4403
rect 154485 4363 154543 4369
rect 154577 4403 154635 4409
rect 154577 4369 154589 4403
rect 154623 4400 154635 4403
rect 164145 4403 164203 4409
rect 164145 4400 164157 4403
rect 154623 4372 164157 4400
rect 154623 4369 154635 4372
rect 154577 4363 154635 4369
rect 164145 4369 164157 4372
rect 164191 4369 164203 4403
rect 164145 4363 164203 4369
rect 215846 4360 215852 4412
rect 215904 4400 215910 4412
rect 247034 4400 247040 4412
rect 215904 4372 247040 4400
rect 215904 4360 215910 4372
rect 247034 4360 247040 4372
rect 247092 4360 247098 4412
rect 251450 4360 251456 4412
rect 251508 4400 251514 4412
rect 255590 4400 255596 4412
rect 251508 4372 255596 4400
rect 251508 4360 251514 4372
rect 255590 4360 255596 4372
rect 255648 4360 255654 4412
rect 258994 4360 259000 4412
rect 259052 4400 259058 4412
rect 263318 4400 263324 4412
rect 259052 4372 263324 4400
rect 259052 4360 259058 4372
rect 263318 4360 263324 4372
rect 263376 4360 263382 4412
rect 263413 4403 263471 4409
rect 263413 4369 263425 4403
rect 263459 4400 263471 4403
rect 264977 4403 265035 4409
rect 263459 4372 264928 4400
rect 263459 4369 263471 4372
rect 263413 4363 263471 4369
rect 176565 4335 176623 4341
rect 176565 4301 176577 4335
rect 176611 4332 176623 4335
rect 180702 4332 180708 4344
rect 176611 4304 180708 4332
rect 176611 4301 176623 4304
rect 176565 4295 176623 4301
rect 180702 4292 180708 4304
rect 180760 4292 180766 4344
rect 215113 4335 215171 4341
rect 215113 4301 215125 4335
rect 215159 4332 215171 4335
rect 215481 4335 215539 4341
rect 215481 4332 215493 4335
rect 215159 4304 215493 4332
rect 215159 4301 215171 4304
rect 215113 4295 215171 4301
rect 215481 4301 215493 4304
rect 215527 4301 215539 4335
rect 215481 4295 215539 4301
rect 219342 4292 219348 4344
rect 219400 4332 219406 4344
rect 239493 4335 239551 4341
rect 219400 4304 239444 4332
rect 219400 4292 219406 4304
rect 215205 4267 215263 4273
rect 215205 4233 215217 4267
rect 215251 4264 215263 4267
rect 215297 4267 215355 4273
rect 215297 4264 215309 4267
rect 215251 4236 215309 4264
rect 215251 4233 215263 4236
rect 215205 4227 215263 4233
rect 215297 4233 215309 4236
rect 215343 4233 215355 4267
rect 215297 4227 215355 4233
rect 222930 4224 222936 4276
rect 222988 4264 222994 4276
rect 239416 4264 239444 4304
rect 239493 4301 239505 4335
rect 239539 4332 239551 4335
rect 249886 4332 249892 4344
rect 239539 4304 249892 4332
rect 239539 4301 239551 4304
rect 239493 4295 239551 4301
rect 249886 4292 249892 4304
rect 249944 4292 249950 4344
rect 252646 4292 252652 4344
rect 252704 4332 252710 4344
rect 255866 4332 255872 4344
rect 252704 4304 255872 4332
rect 252704 4292 252710 4304
rect 255866 4292 255872 4304
rect 255924 4292 255930 4344
rect 259178 4292 259184 4344
rect 259236 4332 259242 4344
rect 264793 4335 264851 4341
rect 264793 4332 264805 4335
rect 259236 4304 264805 4332
rect 259236 4292 259242 4304
rect 264793 4301 264805 4304
rect 264839 4301 264851 4335
rect 264793 4295 264851 4301
rect 248414 4264 248420 4276
rect 222988 4236 239352 4264
rect 239416 4236 248420 4264
rect 222988 4224 222994 4236
rect 128265 4199 128323 4205
rect 128265 4165 128277 4199
rect 128311 4196 128323 4199
rect 128357 4199 128415 4205
rect 128357 4196 128369 4199
rect 128311 4168 128369 4196
rect 128311 4165 128323 4168
rect 128265 4159 128323 4165
rect 128357 4165 128369 4168
rect 128403 4165 128415 4199
rect 128357 4159 128415 4165
rect 147585 4199 147643 4205
rect 147585 4165 147597 4199
rect 147631 4196 147643 4199
rect 157245 4199 157303 4205
rect 157245 4196 157257 4199
rect 147631 4168 157257 4196
rect 147631 4165 147643 4168
rect 147585 4159 147643 4165
rect 157245 4165 157257 4168
rect 157291 4165 157303 4199
rect 157245 4159 157303 4165
rect 176473 4199 176531 4205
rect 176473 4165 176485 4199
rect 176519 4196 176531 4199
rect 180705 4199 180763 4205
rect 180705 4196 180717 4199
rect 176519 4168 180717 4196
rect 176519 4165 176531 4168
rect 176473 4159 176531 4165
rect 180705 4165 180717 4168
rect 180751 4165 180763 4199
rect 180705 4159 180763 4165
rect 180797 4199 180855 4205
rect 180797 4165 180809 4199
rect 180843 4196 180855 4199
rect 190365 4199 190423 4205
rect 190365 4196 190377 4199
rect 180843 4168 190377 4196
rect 180843 4165 180855 4168
rect 180797 4159 180855 4165
rect 190365 4165 190377 4168
rect 190411 4165 190423 4199
rect 190365 4159 190423 4165
rect 200117 4199 200175 4205
rect 200117 4165 200129 4199
rect 200163 4196 200175 4199
rect 205729 4199 205787 4205
rect 205729 4196 205741 4199
rect 200163 4168 205741 4196
rect 200163 4165 200175 4168
rect 200117 4159 200175 4165
rect 205729 4165 205741 4168
rect 205775 4165 205787 4199
rect 205729 4159 205787 4165
rect 215021 4199 215079 4205
rect 215021 4165 215033 4199
rect 215067 4196 215079 4199
rect 215389 4199 215447 4205
rect 215389 4196 215401 4199
rect 215067 4168 215401 4196
rect 215067 4165 215079 4168
rect 215021 4159 215079 4165
rect 215389 4165 215401 4168
rect 215435 4165 215447 4199
rect 215389 4159 215447 4165
rect 220173 4199 220231 4205
rect 220173 4165 220185 4199
rect 220219 4196 220231 4199
rect 224865 4199 224923 4205
rect 224865 4196 224877 4199
rect 220219 4168 224877 4196
rect 220219 4165 220231 4168
rect 220173 4159 220231 4165
rect 224865 4165 224877 4168
rect 224911 4165 224923 4199
rect 224865 4159 224923 4165
rect 226518 4156 226524 4208
rect 226576 4196 226582 4208
rect 239217 4199 239275 4205
rect 239217 4196 239229 4199
rect 226576 4168 239229 4196
rect 226576 4156 226582 4168
rect 239217 4165 239229 4168
rect 239263 4165 239275 4199
rect 239324 4196 239352 4236
rect 248414 4224 248420 4236
rect 248472 4224 248478 4276
rect 249794 4264 249800 4276
rect 248524 4236 249800 4264
rect 248524 4196 248552 4236
rect 249794 4224 249800 4236
rect 249852 4224 249858 4276
rect 253842 4224 253848 4276
rect 253900 4264 253906 4276
rect 255498 4264 255504 4276
rect 253900 4236 255504 4264
rect 253900 4224 253906 4236
rect 255498 4224 255504 4236
rect 255556 4224 255562 4276
rect 264900 4264 264928 4372
rect 264977 4369 264989 4403
rect 265023 4400 265035 4403
rect 281258 4400 281264 4412
rect 265023 4372 281264 4400
rect 265023 4369 265035 4372
rect 264977 4363 265035 4369
rect 281258 4360 281264 4372
rect 281316 4360 281322 4412
rect 307570 4360 307576 4412
rect 307628 4400 307634 4412
rect 501230 4400 501236 4412
rect 307628 4372 501236 4400
rect 307628 4360 307634 4372
rect 501230 4360 501236 4372
rect 501288 4360 501294 4412
rect 265069 4335 265127 4341
rect 265069 4301 265081 4335
rect 265115 4332 265127 4335
rect 265802 4332 265808 4344
rect 265115 4304 265808 4332
rect 265115 4301 265127 4304
rect 265069 4295 265127 4301
rect 265802 4292 265808 4304
rect 265860 4292 265866 4344
rect 267369 4335 267427 4341
rect 267369 4301 267381 4335
rect 267415 4332 267427 4335
rect 277670 4332 277676 4344
rect 267415 4304 277676 4332
rect 267415 4301 267427 4304
rect 267369 4295 267427 4301
rect 277670 4292 277676 4304
rect 277728 4292 277734 4344
rect 292485 4335 292543 4341
rect 292485 4301 292497 4335
rect 292531 4332 292543 4335
rect 292577 4335 292635 4341
rect 292577 4332 292589 4335
rect 292531 4304 292589 4332
rect 292531 4301 292543 4304
rect 292485 4295 292543 4301
rect 292577 4301 292589 4304
rect 292623 4301 292635 4335
rect 292577 4295 292635 4301
rect 307662 4292 307668 4344
rect 307720 4332 307726 4344
rect 497734 4332 497740 4344
rect 307720 4304 497740 4332
rect 307720 4292 307726 4304
rect 497734 4292 497740 4304
rect 497792 4292 497798 4344
rect 266998 4264 267004 4276
rect 264900 4236 267004 4264
rect 266998 4224 267004 4236
rect 267056 4224 267062 4276
rect 268381 4267 268439 4273
rect 268381 4233 268393 4267
rect 268427 4264 268439 4267
rect 274082 4264 274088 4276
rect 268427 4236 274088 4264
rect 268427 4233 268439 4236
rect 268381 4227 268439 4233
rect 274082 4224 274088 4236
rect 274140 4224 274146 4276
rect 282733 4267 282791 4273
rect 282733 4233 282745 4267
rect 282779 4264 282791 4267
rect 292298 4264 292304 4276
rect 282779 4236 292304 4264
rect 282779 4233 282791 4236
rect 282733 4227 282791 4233
rect 292298 4224 292304 4236
rect 292356 4224 292362 4276
rect 292393 4267 292451 4273
rect 292393 4233 292405 4267
rect 292439 4264 292451 4267
rect 292669 4267 292727 4273
rect 292669 4264 292681 4267
rect 292439 4236 292681 4264
rect 292439 4233 292451 4236
rect 292393 4227 292451 4233
rect 292669 4233 292681 4236
rect 292715 4233 292727 4267
rect 292669 4227 292727 4233
rect 306282 4224 306288 4276
rect 306340 4264 306346 4276
rect 494146 4264 494152 4276
rect 306340 4236 494152 4264
rect 306340 4224 306346 4236
rect 494146 4224 494152 4236
rect 494204 4224 494210 4276
rect 239324 4168 248552 4196
rect 239217 4159 239275 4165
rect 249150 4156 249156 4208
rect 249208 4196 249214 4208
rect 254762 4196 254768 4208
rect 249208 4168 254768 4196
rect 249208 4156 249214 4168
rect 254762 4156 254768 4168
rect 254820 4156 254826 4208
rect 259362 4156 259368 4208
rect 259420 4196 259426 4208
rect 264606 4196 264612 4208
rect 259420 4168 264612 4196
rect 259420 4156 259426 4168
rect 264606 4156 264612 4168
rect 264664 4156 264670 4208
rect 264790 4156 264796 4208
rect 264848 4196 264854 4208
rect 270773 4199 270831 4205
rect 270773 4196 270785 4199
rect 264848 4168 270785 4196
rect 264848 4156 264854 4168
rect 270773 4165 270785 4168
rect 270819 4165 270831 4199
rect 270773 4159 270831 4165
rect 271782 4156 271788 4208
rect 271840 4196 271846 4208
rect 326430 4196 326436 4208
rect 271840 4168 326436 4196
rect 271840 4156 271846 4168
rect 326430 4156 326436 4168
rect 326488 4156 326494 4208
rect 326525 4199 326583 4205
rect 326525 4165 326537 4199
rect 326571 4196 326583 4199
rect 330018 4196 330024 4208
rect 326571 4168 330024 4196
rect 326571 4165 326583 4168
rect 326525 4159 326583 4165
rect 330018 4156 330024 4168
rect 330076 4156 330082 4208
rect 36170 4088 36176 4140
rect 36228 4128 36234 4140
rect 37182 4128 37188 4140
rect 36228 4100 37188 4128
rect 36228 4088 36234 4100
rect 37182 4088 37188 4100
rect 37240 4088 37246 4140
rect 37366 4088 37372 4140
rect 37424 4128 37430 4140
rect 38562 4128 38568 4140
rect 37424 4100 38568 4128
rect 37424 4088 37430 4100
rect 38562 4088 38568 4100
rect 38620 4088 38626 4140
rect 42150 4088 42156 4140
rect 42208 4128 42214 4140
rect 42702 4128 42708 4140
rect 42208 4100 42708 4128
rect 42208 4088 42214 4100
rect 42702 4088 42708 4100
rect 42760 4088 42766 4140
rect 44542 4088 44548 4140
rect 44600 4128 44606 4140
rect 45462 4128 45468 4140
rect 44600 4100 45468 4128
rect 44600 4088 44606 4100
rect 45462 4088 45468 4100
rect 45520 4088 45526 4140
rect 55214 4088 55220 4140
rect 55272 4128 55278 4140
rect 56410 4128 56416 4140
rect 55272 4100 56416 4128
rect 55272 4088 55278 4100
rect 56410 4088 56416 4100
rect 56468 4088 56474 4140
rect 58713 4131 58771 4137
rect 58713 4097 58725 4131
rect 58759 4128 58771 4131
rect 334434 4128 334440 4140
rect 58759 4100 334440 4128
rect 58759 4097 58771 4100
rect 58713 4091 58771 4097
rect 334434 4088 334440 4100
rect 334492 4088 334498 4140
rect 46934 4020 46940 4072
rect 46992 4060 46998 4072
rect 332686 4060 332692 4072
rect 46992 4032 332692 4060
rect 46992 4020 46998 4032
rect 332686 4020 332692 4032
rect 332744 4020 332750 4072
rect 45738 3952 45744 4004
rect 45796 3992 45802 4004
rect 332962 3992 332968 4004
rect 45796 3964 332968 3992
rect 45796 3952 45802 3964
rect 332962 3952 332968 3964
rect 333020 3952 333026 4004
rect 39758 3884 39764 3936
rect 39816 3924 39822 3936
rect 331858 3924 331864 3936
rect 39816 3896 331864 3924
rect 39816 3884 39822 3896
rect 331858 3884 331864 3896
rect 331916 3884 331922 3936
rect 38562 3816 38568 3868
rect 38620 3856 38626 3868
rect 55217 3859 55275 3865
rect 55217 3856 55229 3859
rect 38620 3828 55229 3856
rect 38620 3816 38626 3828
rect 55217 3825 55229 3828
rect 55263 3825 55275 3859
rect 55217 3819 55275 3825
rect 64785 3859 64843 3865
rect 64785 3825 64797 3859
rect 64831 3856 64843 3859
rect 168745 3859 168803 3865
rect 168745 3856 168757 3859
rect 64831 3828 168757 3856
rect 64831 3825 64843 3828
rect 64785 3819 64843 3825
rect 168745 3825 168757 3828
rect 168791 3825 168803 3859
rect 168745 3819 168803 3825
rect 168837 3859 168895 3865
rect 168837 3825 168849 3859
rect 168883 3856 168895 3859
rect 171689 3859 171747 3865
rect 171689 3856 171701 3859
rect 168883 3828 171701 3856
rect 168883 3825 168895 3828
rect 168837 3819 168895 3825
rect 171689 3825 171701 3828
rect 171735 3825 171747 3859
rect 171689 3819 171747 3825
rect 171781 3859 171839 3865
rect 171781 3825 171793 3859
rect 171827 3856 171839 3859
rect 180518 3856 180524 3868
rect 171827 3828 180524 3856
rect 171827 3825 171839 3828
rect 171781 3819 171839 3825
rect 180518 3816 180524 3828
rect 180576 3816 180582 3868
rect 180613 3859 180671 3865
rect 180613 3825 180625 3859
rect 180659 3856 180671 3859
rect 215205 3859 215263 3865
rect 215205 3856 215217 3859
rect 180659 3828 215217 3856
rect 180659 3825 180671 3828
rect 180613 3819 180671 3825
rect 215205 3825 215217 3828
rect 215251 3825 215263 3859
rect 215205 3819 215263 3825
rect 215297 3859 215355 3865
rect 215297 3825 215309 3859
rect 215343 3856 215355 3859
rect 263597 3859 263655 3865
rect 263597 3856 263609 3859
rect 215343 3828 263609 3856
rect 215343 3825 215355 3828
rect 215297 3819 215355 3825
rect 263597 3825 263609 3828
rect 263643 3825 263655 3859
rect 263597 3819 263655 3825
rect 263686 3816 263692 3868
rect 263744 3856 263750 3868
rect 282733 3859 282791 3865
rect 282733 3856 282745 3859
rect 263744 3828 282745 3856
rect 263744 3816 263750 3828
rect 282733 3825 282745 3828
rect 282779 3825 282791 3859
rect 282733 3819 282791 3825
rect 282825 3859 282883 3865
rect 282825 3825 282837 3859
rect 282871 3856 282883 3859
rect 292485 3859 292543 3865
rect 292485 3856 292497 3859
rect 282871 3828 292497 3856
rect 282871 3825 282883 3828
rect 282825 3819 282883 3825
rect 292485 3825 292497 3828
rect 292531 3825 292543 3859
rect 292485 3819 292543 3825
rect 292577 3859 292635 3865
rect 292577 3825 292589 3859
rect 292623 3856 292635 3859
rect 303985 3859 304043 3865
rect 303985 3856 303997 3859
rect 292623 3828 303997 3856
rect 292623 3825 292635 3828
rect 292577 3819 292635 3825
rect 303985 3825 303997 3828
rect 304031 3825 304043 3859
rect 303985 3819 304043 3825
rect 304077 3859 304135 3865
rect 304077 3825 304089 3859
rect 304123 3856 304135 3859
rect 306929 3859 306987 3865
rect 306929 3856 306941 3859
rect 304123 3828 306941 3856
rect 304123 3825 304135 3828
rect 304077 3819 304135 3825
rect 306929 3825 306941 3828
rect 306975 3825 306987 3859
rect 306929 3819 306987 3825
rect 307021 3859 307079 3865
rect 307021 3825 307033 3859
rect 307067 3856 307079 3859
rect 316681 3859 316739 3865
rect 316681 3856 316693 3859
rect 307067 3828 316693 3856
rect 307067 3825 307079 3828
rect 307021 3819 307079 3825
rect 316681 3825 316693 3828
rect 316727 3825 316739 3859
rect 316681 3819 316739 3825
rect 316773 3859 316831 3865
rect 316773 3825 316785 3859
rect 316819 3856 316831 3859
rect 331674 3856 331680 3868
rect 316819 3828 331680 3856
rect 316819 3825 316831 3828
rect 316773 3819 316831 3825
rect 331674 3816 331680 3828
rect 331732 3816 331738 3868
rect 32674 3748 32680 3800
rect 32732 3788 32738 3800
rect 329926 3788 329932 3800
rect 32732 3760 329932 3788
rect 32732 3748 32738 3760
rect 329926 3748 329932 3760
rect 329984 3748 329990 3800
rect 31478 3680 31484 3732
rect 31536 3720 31542 3732
rect 55217 3723 55275 3729
rect 55217 3720 55229 3723
rect 31536 3692 55229 3720
rect 31536 3680 31542 3692
rect 55217 3689 55229 3692
rect 55263 3689 55275 3723
rect 55217 3683 55275 3689
rect 64785 3723 64843 3729
rect 64785 3689 64797 3723
rect 64831 3720 64843 3723
rect 171965 3723 172023 3729
rect 64831 3692 171916 3720
rect 64831 3689 64843 3692
rect 64785 3683 64843 3689
rect 27890 3612 27896 3664
rect 27948 3652 27954 3664
rect 34609 3655 34667 3661
rect 27948 3624 34560 3652
rect 27948 3612 27954 3624
rect 12434 3544 12440 3596
rect 12492 3584 12498 3596
rect 13630 3584 13636 3596
rect 12492 3556 13636 3584
rect 12492 3544 12498 3556
rect 13630 3544 13636 3556
rect 13688 3544 13694 3596
rect 26694 3544 26700 3596
rect 26752 3584 26758 3596
rect 27522 3584 27528 3596
rect 26752 3556 27528 3584
rect 26752 3544 26758 3556
rect 27522 3544 27528 3556
rect 27580 3544 27586 3596
rect 33870 3544 33876 3596
rect 33928 3584 33934 3596
rect 34422 3584 34428 3596
rect 33928 3556 34428 3584
rect 33928 3544 33934 3556
rect 34422 3544 34428 3556
rect 34480 3544 34486 3596
rect 34532 3584 34560 3624
rect 34609 3621 34621 3655
rect 34655 3652 34667 3655
rect 64877 3655 64935 3661
rect 64877 3652 64889 3655
rect 34655 3624 55352 3652
rect 34655 3621 34667 3624
rect 34609 3615 34667 3621
rect 55217 3587 55275 3593
rect 55217 3584 55229 3587
rect 34532 3556 55229 3584
rect 55217 3553 55229 3556
rect 55263 3553 55275 3587
rect 55324 3584 55352 3624
rect 64708 3624 64889 3652
rect 64708 3584 64736 3624
rect 64877 3621 64889 3624
rect 64923 3621 64935 3655
rect 64877 3615 64935 3621
rect 74445 3655 74503 3661
rect 74445 3621 74457 3655
rect 74491 3652 74503 3655
rect 84197 3655 84255 3661
rect 84197 3652 84209 3655
rect 74491 3624 84209 3652
rect 74491 3621 74503 3624
rect 74445 3615 74503 3621
rect 84197 3621 84209 3624
rect 84243 3621 84255 3655
rect 84197 3615 84255 3621
rect 93302 3612 93308 3664
rect 93360 3652 93366 3664
rect 93762 3652 93768 3664
rect 93360 3624 93768 3652
rect 93360 3612 93366 3624
rect 93762 3612 93768 3624
rect 93820 3612 93826 3664
rect 94498 3612 94504 3664
rect 94556 3652 94562 3664
rect 95142 3652 95148 3664
rect 94556 3624 95148 3652
rect 94556 3612 94562 3624
rect 95142 3612 95148 3624
rect 95200 3612 95206 3664
rect 95694 3612 95700 3664
rect 95752 3652 95758 3664
rect 96522 3652 96528 3664
rect 95752 3624 96528 3652
rect 95752 3612 95758 3624
rect 96522 3612 96528 3624
rect 96580 3612 96586 3664
rect 98086 3612 98092 3664
rect 98144 3652 98150 3664
rect 99190 3652 99196 3664
rect 98144 3624 99196 3652
rect 98144 3612 98150 3624
rect 99190 3612 99196 3624
rect 99248 3612 99254 3664
rect 99285 3655 99343 3661
rect 99285 3621 99297 3655
rect 99331 3652 99343 3655
rect 101493 3655 101551 3661
rect 101493 3652 101505 3655
rect 99331 3624 101505 3652
rect 99331 3621 99343 3624
rect 99285 3615 99343 3621
rect 101493 3621 101505 3624
rect 101539 3621 101551 3655
rect 101493 3615 101551 3621
rect 101582 3612 101588 3664
rect 101640 3652 101646 3664
rect 102042 3652 102048 3664
rect 101640 3624 102048 3652
rect 101640 3612 101646 3624
rect 102042 3612 102048 3624
rect 102100 3612 102106 3664
rect 102778 3612 102784 3664
rect 102836 3652 102842 3664
rect 103422 3652 103428 3664
rect 102836 3624 103428 3652
rect 102836 3612 102842 3624
rect 103422 3612 103428 3624
rect 103480 3612 103486 3664
rect 105170 3612 105176 3664
rect 105228 3652 105234 3664
rect 106182 3652 106188 3664
rect 105228 3624 106188 3652
rect 105228 3612 105234 3624
rect 106182 3612 106188 3624
rect 106240 3612 106246 3664
rect 112346 3612 112352 3664
rect 112404 3652 112410 3664
rect 113082 3652 113088 3664
rect 112404 3624 113088 3652
rect 112404 3612 112410 3624
rect 113082 3612 113088 3624
rect 113140 3612 113146 3664
rect 114738 3612 114744 3664
rect 114796 3652 114802 3664
rect 115842 3652 115848 3664
rect 114796 3624 115848 3652
rect 114796 3612 114802 3624
rect 115842 3612 115848 3624
rect 115900 3612 115906 3664
rect 115934 3612 115940 3664
rect 115992 3652 115998 3664
rect 117222 3652 117228 3664
rect 115992 3624 117228 3652
rect 115992 3612 115998 3624
rect 117222 3612 117228 3624
rect 117280 3612 117286 3664
rect 117317 3655 117375 3661
rect 117317 3621 117329 3655
rect 117363 3652 117375 3655
rect 119341 3655 119399 3661
rect 119341 3652 119353 3655
rect 117363 3624 119353 3652
rect 117363 3621 117375 3624
rect 117317 3615 117375 3621
rect 119341 3621 119353 3624
rect 119387 3621 119399 3655
rect 119341 3615 119399 3621
rect 119430 3612 119436 3664
rect 119488 3652 119494 3664
rect 119982 3652 119988 3664
rect 119488 3624 119988 3652
rect 119488 3612 119494 3624
rect 119982 3612 119988 3624
rect 120040 3612 120046 3664
rect 121822 3612 121828 3664
rect 121880 3652 121886 3664
rect 122742 3652 122748 3664
rect 121880 3624 122748 3652
rect 121880 3612 121886 3624
rect 122742 3612 122748 3624
rect 122800 3612 122806 3664
rect 123018 3612 123024 3664
rect 123076 3652 123082 3664
rect 124122 3652 124128 3664
rect 123076 3624 124128 3652
rect 123076 3612 123082 3624
rect 124122 3612 124128 3624
rect 124180 3612 124186 3664
rect 124217 3655 124275 3661
rect 124217 3621 124229 3655
rect 124263 3652 124275 3655
rect 128265 3655 128323 3661
rect 128265 3652 128277 3655
rect 124263 3624 128277 3652
rect 124263 3621 124275 3624
rect 124217 3615 124275 3621
rect 128265 3621 128277 3624
rect 128311 3621 128323 3655
rect 128265 3615 128323 3621
rect 128357 3655 128415 3661
rect 128357 3621 128369 3655
rect 128403 3652 128415 3655
rect 147585 3655 147643 3661
rect 147585 3652 147597 3655
rect 128403 3624 147597 3652
rect 128403 3621 128415 3624
rect 128357 3615 128415 3621
rect 147585 3621 147597 3624
rect 147631 3621 147643 3655
rect 147585 3615 147643 3621
rect 157245 3655 157303 3661
rect 157245 3621 157257 3655
rect 157291 3652 157303 3655
rect 171781 3655 171839 3661
rect 171781 3652 171793 3655
rect 157291 3624 171793 3652
rect 157291 3621 157303 3624
rect 157245 3615 157303 3621
rect 171781 3621 171793 3624
rect 171827 3621 171839 3655
rect 171888 3652 171916 3692
rect 171965 3689 171977 3723
rect 172011 3720 172023 3723
rect 180521 3723 180579 3729
rect 180521 3720 180533 3723
rect 172011 3692 180533 3720
rect 172011 3689 172023 3692
rect 171965 3683 172023 3689
rect 180521 3689 180533 3692
rect 180567 3689 180579 3723
rect 180521 3683 180579 3689
rect 180610 3680 180616 3732
rect 180668 3680 180674 3732
rect 180702 3680 180708 3732
rect 180760 3720 180766 3732
rect 205729 3723 205787 3729
rect 180760 3692 205680 3720
rect 180760 3680 180766 3692
rect 176565 3655 176623 3661
rect 176565 3652 176577 3655
rect 171888 3624 176577 3652
rect 171781 3615 171839 3621
rect 176565 3621 176577 3624
rect 176611 3621 176623 3655
rect 180628 3652 180656 3680
rect 180797 3655 180855 3661
rect 180797 3652 180809 3655
rect 180628 3624 180809 3652
rect 176565 3615 176623 3621
rect 180797 3621 180809 3624
rect 180843 3621 180855 3655
rect 180797 3615 180855 3621
rect 190365 3655 190423 3661
rect 190365 3621 190377 3655
rect 190411 3652 190423 3655
rect 200117 3655 200175 3661
rect 200117 3652 200129 3655
rect 190411 3624 200129 3652
rect 190411 3621 190423 3624
rect 190365 3615 190423 3621
rect 200117 3621 200129 3624
rect 200163 3621 200175 3655
rect 205652 3652 205680 3692
rect 205729 3689 205741 3723
rect 205775 3720 205787 3723
rect 215389 3723 215447 3729
rect 205775 3692 215340 3720
rect 205775 3689 205787 3692
rect 205729 3683 205787 3689
rect 215113 3655 215171 3661
rect 215113 3652 215125 3655
rect 205652 3624 215125 3652
rect 200117 3615 200175 3621
rect 215113 3621 215125 3624
rect 215159 3621 215171 3655
rect 215312 3652 215340 3692
rect 215389 3689 215401 3723
rect 215435 3720 215447 3723
rect 220173 3723 220231 3729
rect 220173 3720 220185 3723
rect 215435 3692 220185 3720
rect 215435 3689 215447 3692
rect 215389 3683 215447 3689
rect 220173 3689 220185 3692
rect 220219 3689 220231 3723
rect 220173 3683 220231 3689
rect 220265 3723 220323 3729
rect 220265 3689 220277 3723
rect 220311 3720 220323 3723
rect 273070 3720 273076 3732
rect 220311 3692 273076 3720
rect 220311 3689 220323 3692
rect 220265 3683 220323 3689
rect 273070 3680 273076 3692
rect 273128 3680 273134 3732
rect 273346 3680 273352 3732
rect 273404 3720 273410 3732
rect 292390 3720 292396 3732
rect 273404 3692 292396 3720
rect 273404 3680 273410 3692
rect 292390 3680 292396 3692
rect 292448 3680 292454 3732
rect 292482 3680 292488 3732
rect 292540 3720 292546 3732
rect 292540 3692 292620 3720
rect 292540 3680 292546 3692
rect 224770 3652 224776 3664
rect 215312 3624 224776 3652
rect 215113 3615 215171 3621
rect 224770 3612 224776 3624
rect 224828 3612 224834 3664
rect 224954 3612 224960 3664
rect 225012 3652 225018 3664
rect 263410 3652 263416 3664
rect 225012 3624 263416 3652
rect 225012 3612 225018 3624
rect 263410 3612 263416 3624
rect 263468 3612 263474 3664
rect 270497 3655 270555 3661
rect 270497 3652 270509 3655
rect 263520 3624 270509 3652
rect 55324 3556 64736 3584
rect 64785 3587 64843 3593
rect 55217 3547 55275 3553
rect 64785 3553 64797 3587
rect 64831 3584 64843 3587
rect 168653 3587 168711 3593
rect 168653 3584 168665 3587
rect 64831 3556 168665 3584
rect 64831 3553 64843 3556
rect 64785 3547 64843 3553
rect 168653 3553 168665 3556
rect 168699 3553 168711 3587
rect 168653 3547 168711 3553
rect 168745 3587 168803 3593
rect 168745 3553 168757 3587
rect 168791 3584 168803 3587
rect 180613 3587 180671 3593
rect 180613 3584 180625 3587
rect 168791 3556 180625 3584
rect 168791 3553 168803 3556
rect 168745 3547 168803 3553
rect 180613 3553 180625 3556
rect 180659 3553 180671 3587
rect 180613 3547 180671 3553
rect 180705 3587 180763 3593
rect 180705 3553 180717 3587
rect 180751 3584 180763 3587
rect 208029 3587 208087 3593
rect 208029 3584 208041 3587
rect 180751 3556 208041 3584
rect 180751 3553 180763 3556
rect 180705 3547 180763 3553
rect 208029 3553 208041 3556
rect 208075 3553 208087 3587
rect 208029 3547 208087 3553
rect 208121 3587 208179 3593
rect 208121 3553 208133 3587
rect 208167 3584 208179 3587
rect 220081 3587 220139 3593
rect 220081 3584 220093 3587
rect 208167 3556 220093 3584
rect 208167 3553 208179 3556
rect 208121 3547 208179 3553
rect 220081 3553 220093 3556
rect 220127 3553 220139 3587
rect 220081 3547 220139 3553
rect 224865 3587 224923 3593
rect 224865 3553 224877 3587
rect 224911 3584 224923 3587
rect 263520 3584 263548 3624
rect 270497 3621 270509 3624
rect 270543 3621 270555 3655
rect 292592 3652 292620 3692
rect 292666 3680 292672 3732
rect 292724 3720 292730 3732
rect 303801 3723 303859 3729
rect 303801 3720 303813 3723
rect 292724 3692 303813 3720
rect 292724 3680 292730 3692
rect 303801 3689 303813 3692
rect 303847 3689 303859 3723
rect 303801 3683 303859 3689
rect 303893 3723 303951 3729
rect 303893 3689 303905 3723
rect 303939 3720 303951 3723
rect 306837 3723 306895 3729
rect 306837 3720 306849 3723
rect 303939 3692 306849 3720
rect 303939 3689 303951 3692
rect 303893 3683 303951 3689
rect 306837 3689 306849 3692
rect 306883 3689 306895 3723
rect 306837 3683 306895 3689
rect 306929 3723 306987 3729
rect 306929 3689 306941 3723
rect 306975 3720 306987 3723
rect 313737 3723 313795 3729
rect 313737 3720 313749 3723
rect 306975 3692 313749 3720
rect 306975 3689 306987 3692
rect 306929 3683 306987 3689
rect 313737 3689 313749 3692
rect 313783 3689 313795 3723
rect 313737 3683 313795 3689
rect 313844 3692 316908 3720
rect 307021 3655 307079 3661
rect 307021 3652 307033 3655
rect 292592 3624 307033 3652
rect 270497 3615 270555 3621
rect 307021 3621 307033 3624
rect 307067 3621 307079 3655
rect 307021 3615 307079 3621
rect 307113 3655 307171 3661
rect 307113 3621 307125 3655
rect 307159 3652 307171 3655
rect 311802 3652 311808 3664
rect 307159 3624 311808 3652
rect 307159 3621 307171 3624
rect 307113 3615 307171 3621
rect 311802 3612 311808 3624
rect 311860 3612 311866 3664
rect 313645 3655 313703 3661
rect 313645 3621 313657 3655
rect 313691 3652 313703 3655
rect 313844 3652 313872 3692
rect 313691 3624 313872 3652
rect 313691 3621 313703 3624
rect 313645 3615 313703 3621
rect 313918 3612 313924 3664
rect 313976 3652 313982 3664
rect 316586 3652 316592 3664
rect 313976 3624 316592 3652
rect 313976 3612 313982 3624
rect 316586 3612 316592 3624
rect 316644 3612 316650 3664
rect 224911 3556 263548 3584
rect 263689 3587 263747 3593
rect 224911 3553 224923 3556
rect 224865 3547 224923 3553
rect 263689 3553 263701 3587
rect 263735 3584 263747 3587
rect 265989 3587 266047 3593
rect 265989 3584 266001 3587
rect 263735 3556 266001 3584
rect 263735 3553 263747 3556
rect 263689 3547 263747 3553
rect 265989 3553 266001 3556
rect 266035 3553 266047 3587
rect 265989 3547 266047 3553
rect 266081 3587 266139 3593
rect 266081 3553 266093 3587
rect 266127 3584 266139 3587
rect 278041 3587 278099 3593
rect 278041 3584 278053 3587
rect 266127 3556 278053 3584
rect 266127 3553 266139 3556
rect 266081 3547 266139 3553
rect 278041 3553 278053 3556
rect 278087 3553 278099 3587
rect 278041 3547 278099 3553
rect 278133 3587 278191 3593
rect 278133 3553 278145 3587
rect 278179 3584 278191 3587
rect 282733 3587 282791 3593
rect 282733 3584 282745 3587
rect 278179 3556 282745 3584
rect 278179 3553 278191 3556
rect 278133 3547 278191 3553
rect 282733 3553 282745 3556
rect 282779 3553 282791 3587
rect 282733 3547 282791 3553
rect 282822 3544 282828 3596
rect 282880 3584 282886 3596
rect 285309 3587 285367 3593
rect 285309 3584 285321 3587
rect 282880 3556 285321 3584
rect 282880 3544 282886 3556
rect 285309 3553 285321 3556
rect 285355 3553 285367 3587
rect 285309 3547 285367 3553
rect 285401 3587 285459 3593
rect 285401 3553 285413 3587
rect 285447 3584 285459 3587
rect 297361 3587 297419 3593
rect 297361 3584 297373 3587
rect 285447 3556 297373 3584
rect 285447 3553 285459 3556
rect 285401 3547 285459 3553
rect 297361 3553 297373 3556
rect 297407 3553 297419 3587
rect 297361 3547 297419 3553
rect 297453 3587 297511 3593
rect 297453 3553 297465 3587
rect 297499 3584 297511 3587
rect 303893 3587 303951 3593
rect 303893 3584 303905 3587
rect 297499 3556 303905 3584
rect 297499 3553 297511 3556
rect 297453 3547 297511 3553
rect 303893 3553 303905 3556
rect 303939 3553 303951 3587
rect 303893 3547 303951 3553
rect 303985 3587 304043 3593
rect 303985 3553 303997 3587
rect 304031 3584 304043 3587
rect 316773 3587 316831 3593
rect 316773 3584 316785 3587
rect 304031 3556 316785 3584
rect 304031 3553 304043 3556
rect 303985 3547 304043 3553
rect 316773 3553 316785 3556
rect 316819 3553 316831 3587
rect 316880 3584 316908 3692
rect 316954 3680 316960 3732
rect 317012 3720 317018 3732
rect 324866 3720 324872 3732
rect 317012 3692 324872 3720
rect 317012 3680 317018 3692
rect 324866 3680 324872 3692
rect 324924 3680 324930 3732
rect 324961 3723 325019 3729
rect 324961 3689 324973 3723
rect 325007 3720 325019 3723
rect 328914 3720 328920 3732
rect 325007 3692 328920 3720
rect 325007 3689 325019 3692
rect 324961 3683 325019 3689
rect 328914 3680 328920 3692
rect 328972 3680 328978 3732
rect 317049 3655 317107 3661
rect 317049 3621 317061 3655
rect 317095 3652 317107 3655
rect 326249 3655 326307 3661
rect 326249 3652 326261 3655
rect 317095 3624 326261 3652
rect 317095 3621 317107 3624
rect 317049 3615 317107 3621
rect 326249 3621 326261 3624
rect 326295 3621 326307 3655
rect 326249 3615 326307 3621
rect 326617 3655 326675 3661
rect 326617 3621 326629 3655
rect 326663 3652 326675 3655
rect 337194 3652 337200 3664
rect 326663 3624 337200 3652
rect 326663 3621 326675 3624
rect 326617 3615 326675 3621
rect 337194 3612 337200 3624
rect 337252 3612 337258 3664
rect 433426 3612 433432 3664
rect 433484 3652 433490 3664
rect 434622 3652 434628 3664
rect 433484 3624 434628 3652
rect 433484 3612 433490 3624
rect 434622 3612 434628 3624
rect 434680 3612 434686 3664
rect 477494 3612 477500 3664
rect 477552 3652 477558 3664
rect 478690 3652 478696 3664
rect 477552 3624 478696 3652
rect 477552 3612 477558 3624
rect 478690 3612 478696 3624
rect 478748 3612 478754 3664
rect 485774 3612 485780 3664
rect 485832 3652 485838 3664
rect 486970 3652 486976 3664
rect 485832 3624 486976 3652
rect 485832 3612 485838 3624
rect 486970 3612 486976 3624
rect 487028 3612 487034 3664
rect 316880 3556 325372 3584
rect 316773 3547 316831 3553
rect 566 3476 572 3528
rect 624 3516 630 3528
rect 1302 3516 1308 3528
rect 624 3488 1308 3516
rect 624 3476 630 3488
rect 1302 3476 1308 3488
rect 1360 3476 1366 3528
rect 1670 3476 1676 3528
rect 1728 3516 1734 3528
rect 2682 3516 2688 3528
rect 1728 3488 2688 3516
rect 1728 3476 1734 3488
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 3970 3516 3976 3528
rect 2924 3488 3976 3516
rect 2924 3476 2930 3488
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 8202 3516 8208 3528
rect 7708 3488 8208 3516
rect 7708 3476 7714 3488
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 8846 3476 8852 3528
rect 8904 3516 8910 3528
rect 9582 3516 9588 3528
rect 8904 3488 9588 3516
rect 8904 3476 8910 3488
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 10042 3476 10048 3528
rect 10100 3516 10106 3528
rect 10962 3516 10968 3528
rect 10100 3488 10968 3516
rect 10100 3476 10106 3488
rect 10962 3476 10968 3488
rect 11020 3476 11026 3528
rect 11238 3476 11244 3528
rect 11296 3516 11302 3528
rect 12342 3516 12348 3528
rect 11296 3488 12348 3516
rect 11296 3476 11302 3488
rect 12342 3476 12348 3488
rect 12400 3476 12406 3528
rect 17218 3476 17224 3528
rect 17276 3516 17282 3528
rect 17862 3516 17868 3528
rect 17276 3488 17868 3516
rect 17276 3476 17282 3488
rect 17862 3476 17868 3488
rect 17920 3476 17926 3528
rect 25498 3476 25504 3528
rect 25556 3516 25562 3528
rect 324961 3519 325019 3525
rect 324961 3516 324973 3519
rect 25556 3488 324973 3516
rect 25556 3476 25562 3488
rect 324961 3485 324973 3488
rect 325007 3485 325019 3519
rect 325344 3516 325372 3556
rect 327074 3544 327080 3596
rect 327132 3584 327138 3596
rect 566734 3584 566740 3596
rect 327132 3556 566740 3584
rect 327132 3544 327138 3556
rect 566734 3544 566740 3556
rect 566792 3544 566798 3596
rect 325344 3488 328040 3516
rect 324961 3479 325019 3485
rect 19518 3408 19524 3460
rect 19576 3448 19582 3460
rect 327810 3448 327816 3460
rect 19576 3420 327816 3448
rect 19576 3408 19582 3420
rect 327810 3408 327816 3420
rect 327868 3408 327874 3460
rect 29086 3340 29092 3392
rect 29144 3380 29150 3392
rect 34609 3383 34667 3389
rect 34609 3380 34621 3383
rect 29144 3352 34621 3380
rect 29144 3340 29150 3352
rect 34609 3349 34621 3352
rect 34655 3349 34667 3383
rect 34609 3343 34667 3349
rect 51626 3340 51632 3392
rect 51684 3380 51690 3392
rect 52362 3380 52368 3392
rect 51684 3352 52368 3380
rect 51684 3340 51690 3352
rect 52362 3340 52368 3352
rect 52420 3340 52426 3392
rect 52822 3340 52828 3392
rect 52880 3380 52886 3392
rect 53742 3380 53748 3392
rect 52880 3352 53748 3380
rect 52880 3340 52886 3352
rect 53742 3340 53748 3352
rect 53800 3340 53806 3392
rect 58713 3383 58771 3389
rect 58713 3380 58725 3383
rect 53852 3352 58725 3380
rect 50522 3272 50528 3324
rect 50580 3312 50586 3324
rect 53852 3312 53880 3352
rect 58713 3349 58725 3352
rect 58759 3349 58771 3383
rect 58713 3343 58771 3349
rect 58802 3340 58808 3392
rect 58860 3380 58866 3392
rect 59262 3380 59268 3392
rect 58860 3352 59268 3380
rect 58860 3340 58866 3352
rect 59262 3340 59268 3352
rect 59320 3340 59326 3392
rect 59998 3340 60004 3392
rect 60056 3380 60062 3392
rect 60642 3380 60648 3392
rect 60056 3352 60648 3380
rect 60056 3340 60062 3352
rect 60642 3340 60648 3352
rect 60700 3340 60706 3392
rect 61194 3340 61200 3392
rect 61252 3380 61258 3392
rect 62022 3380 62028 3392
rect 61252 3352 62028 3380
rect 61252 3340 61258 3352
rect 62022 3340 62028 3352
rect 62080 3340 62086 3392
rect 62390 3340 62396 3392
rect 62448 3380 62454 3392
rect 63402 3380 63408 3392
rect 62448 3352 63408 3380
rect 62448 3340 62454 3352
rect 63402 3340 63408 3352
rect 63460 3340 63466 3392
rect 63586 3340 63592 3392
rect 63644 3380 63650 3392
rect 64782 3380 64788 3392
rect 63644 3352 64788 3380
rect 63644 3340 63650 3352
rect 64782 3340 64788 3352
rect 64840 3340 64846 3392
rect 68278 3340 68284 3392
rect 68336 3380 68342 3392
rect 68922 3380 68928 3392
rect 68336 3352 68928 3380
rect 68336 3340 68342 3352
rect 68922 3340 68928 3352
rect 68980 3340 68986 3392
rect 69474 3340 69480 3392
rect 69532 3380 69538 3392
rect 70302 3380 70308 3392
rect 69532 3352 70308 3380
rect 69532 3340 69538 3352
rect 70302 3340 70308 3352
rect 70360 3340 70366 3392
rect 70670 3340 70676 3392
rect 70728 3380 70734 3392
rect 71682 3380 71688 3392
rect 70728 3352 71688 3380
rect 70728 3340 70734 3352
rect 71682 3340 71688 3352
rect 71740 3340 71746 3392
rect 171781 3383 171839 3389
rect 171781 3380 171793 3383
rect 71792 3352 171793 3380
rect 50580 3284 53880 3312
rect 50580 3272 50586 3284
rect 54018 3272 54024 3324
rect 54076 3312 54082 3324
rect 55122 3312 55128 3324
rect 54076 3284 55128 3312
rect 54076 3272 54082 3284
rect 55122 3272 55128 3284
rect 55180 3272 55186 3324
rect 55217 3315 55275 3321
rect 55217 3281 55229 3315
rect 55263 3312 55275 3315
rect 64693 3315 64751 3321
rect 64693 3312 64705 3315
rect 55263 3284 64705 3312
rect 55263 3281 55275 3284
rect 55217 3275 55275 3281
rect 64693 3281 64705 3284
rect 64739 3281 64751 3315
rect 64693 3275 64751 3281
rect 43346 3204 43352 3256
rect 43404 3244 43410 3256
rect 44082 3244 44088 3256
rect 43404 3216 44088 3244
rect 43404 3204 43410 3216
rect 44082 3204 44088 3216
rect 44140 3204 44146 3256
rect 55309 3247 55367 3253
rect 55309 3213 55321 3247
rect 55355 3244 55367 3247
rect 64601 3247 64659 3253
rect 64601 3244 64613 3247
rect 55355 3216 64613 3244
rect 55355 3213 55367 3216
rect 55309 3207 55367 3213
rect 64601 3213 64613 3216
rect 64647 3213 64659 3247
rect 64601 3207 64659 3213
rect 64782 3204 64788 3256
rect 64840 3244 64846 3256
rect 71792 3244 71820 3352
rect 171781 3349 171793 3352
rect 171827 3349 171839 3383
rect 171781 3343 171839 3349
rect 171873 3383 171931 3389
rect 171873 3349 171885 3383
rect 171919 3380 171931 3383
rect 176473 3383 176531 3389
rect 176473 3380 176485 3383
rect 171919 3352 176485 3380
rect 171919 3349 171931 3352
rect 171873 3343 171931 3349
rect 176473 3349 176485 3352
rect 176519 3349 176531 3383
rect 176473 3343 176531 3349
rect 180705 3383 180763 3389
rect 180705 3349 180717 3383
rect 180751 3380 180763 3383
rect 208121 3383 208179 3389
rect 208121 3380 208133 3383
rect 180751 3352 208133 3380
rect 180751 3349 180763 3352
rect 180705 3343 180763 3349
rect 208121 3349 208133 3352
rect 208167 3349 208179 3383
rect 208121 3343 208179 3349
rect 208213 3383 208271 3389
rect 208213 3349 208225 3383
rect 208259 3380 208271 3383
rect 215021 3383 215079 3389
rect 215021 3380 215033 3383
rect 208259 3352 215033 3380
rect 208259 3349 208271 3352
rect 208213 3343 208271 3349
rect 215021 3349 215033 3352
rect 215067 3349 215079 3383
rect 215021 3343 215079 3349
rect 215481 3383 215539 3389
rect 215481 3349 215493 3383
rect 215527 3380 215539 3383
rect 219989 3383 220047 3389
rect 219989 3380 220001 3383
rect 215527 3352 220001 3380
rect 215527 3349 215539 3352
rect 215481 3343 215539 3349
rect 219989 3349 220001 3352
rect 220035 3349 220047 3383
rect 219989 3343 220047 3349
rect 220081 3383 220139 3389
rect 220081 3349 220093 3383
rect 220127 3380 220139 3383
rect 266081 3383 266139 3389
rect 266081 3380 266093 3383
rect 220127 3352 266093 3380
rect 220127 3349 220139 3352
rect 220081 3343 220139 3349
rect 266081 3349 266093 3352
rect 266127 3349 266139 3383
rect 266081 3343 266139 3349
rect 266173 3383 266231 3389
rect 266173 3349 266185 3383
rect 266219 3380 266231 3383
rect 267737 3383 267795 3389
rect 267737 3380 267749 3383
rect 266219 3352 267749 3380
rect 266219 3349 266231 3352
rect 266173 3343 266231 3349
rect 267737 3349 267749 3352
rect 267783 3349 267795 3383
rect 267737 3343 267795 3349
rect 270497 3383 270555 3389
rect 270497 3349 270509 3383
rect 270543 3380 270555 3383
rect 275186 3380 275192 3392
rect 270543 3352 275192 3380
rect 270543 3349 270555 3352
rect 270497 3343 270555 3349
rect 275186 3340 275192 3352
rect 275244 3340 275250 3392
rect 277305 3383 277363 3389
rect 277305 3349 277317 3383
rect 277351 3380 277363 3383
rect 277949 3383 278007 3389
rect 277949 3380 277961 3383
rect 277351 3352 277961 3380
rect 277351 3349 277363 3352
rect 277305 3343 277363 3349
rect 277949 3349 277961 3352
rect 277995 3349 278007 3383
rect 277949 3343 278007 3349
rect 278041 3383 278099 3389
rect 278041 3349 278053 3383
rect 278087 3380 278099 3383
rect 285401 3383 285459 3389
rect 285401 3380 285413 3383
rect 278087 3352 285413 3380
rect 278087 3349 278099 3352
rect 278041 3343 278099 3349
rect 285401 3349 285413 3352
rect 285447 3349 285459 3383
rect 285401 3343 285459 3349
rect 285493 3383 285551 3389
rect 285493 3349 285505 3383
rect 285539 3380 285551 3383
rect 292393 3383 292451 3389
rect 292393 3380 292405 3383
rect 285539 3352 292405 3380
rect 285539 3349 285551 3352
rect 285493 3343 285551 3349
rect 292393 3349 292405 3352
rect 292439 3349 292451 3383
rect 292393 3343 292451 3349
rect 292669 3383 292727 3389
rect 292669 3349 292681 3383
rect 292715 3380 292727 3383
rect 297269 3383 297327 3389
rect 297269 3380 297281 3383
rect 292715 3352 297281 3380
rect 292715 3349 292727 3352
rect 292669 3343 292727 3349
rect 297269 3349 297281 3352
rect 297315 3349 297327 3383
rect 297269 3343 297327 3349
rect 297361 3383 297419 3389
rect 297361 3349 297373 3383
rect 297407 3380 297419 3383
rect 306929 3383 306987 3389
rect 306929 3380 306941 3383
rect 297407 3352 306941 3380
rect 297407 3349 297419 3352
rect 297361 3343 297419 3349
rect 306929 3349 306941 3352
rect 306975 3349 306987 3383
rect 306929 3343 306987 3349
rect 307021 3383 307079 3389
rect 307021 3349 307033 3383
rect 307067 3380 307079 3383
rect 313645 3383 313703 3389
rect 313645 3380 313657 3383
rect 307067 3352 313657 3380
rect 307067 3349 307079 3352
rect 307021 3343 307079 3349
rect 313645 3349 313657 3352
rect 313691 3349 313703 3383
rect 313645 3343 313703 3349
rect 313737 3383 313795 3389
rect 313737 3349 313749 3383
rect 313783 3380 313795 3383
rect 326617 3383 326675 3389
rect 326617 3380 326629 3383
rect 313783 3352 326629 3380
rect 313783 3349 313795 3352
rect 313737 3343 313795 3349
rect 326617 3349 326629 3352
rect 326663 3349 326675 3383
rect 328012 3380 328040 3488
rect 328638 3476 328644 3528
rect 328696 3516 328702 3528
rect 571426 3516 571432 3528
rect 328696 3488 571432 3516
rect 328696 3476 328702 3488
rect 571426 3476 571432 3488
rect 571484 3476 571490 3528
rect 580994 3476 581000 3528
rect 581052 3516 581058 3528
rect 582190 3516 582196 3528
rect 581052 3488 582196 3516
rect 581052 3476 581058 3488
rect 582190 3476 582196 3488
rect 582248 3476 582254 3528
rect 328454 3408 328460 3460
rect 328512 3448 328518 3460
rect 573818 3448 573824 3460
rect 328512 3420 573824 3448
rect 328512 3408 328518 3420
rect 573818 3408 573824 3420
rect 573876 3408 573882 3460
rect 329190 3380 329196 3392
rect 328012 3352 329196 3380
rect 326617 3343 326675 3349
rect 329190 3340 329196 3352
rect 329248 3340 329254 3392
rect 373994 3340 374000 3392
rect 374052 3380 374058 3392
rect 375190 3380 375196 3392
rect 374052 3352 375196 3380
rect 374052 3340 374058 3352
rect 375190 3340 375196 3352
rect 375248 3340 375254 3392
rect 390554 3340 390560 3392
rect 390612 3380 390618 3392
rect 391842 3380 391848 3392
rect 390612 3352 391848 3380
rect 390612 3340 390618 3352
rect 391842 3340 391848 3352
rect 391900 3340 391906 3392
rect 408494 3340 408500 3392
rect 408552 3380 408558 3392
rect 409690 3380 409696 3392
rect 408552 3352 409696 3380
rect 408552 3340 408558 3352
rect 409690 3340 409696 3352
rect 409748 3340 409754 3392
rect 416774 3340 416780 3392
rect 416832 3380 416838 3392
rect 417970 3380 417976 3392
rect 416832 3352 417976 3380
rect 416832 3340 416838 3352
rect 417970 3340 417976 3352
rect 418028 3340 418034 3392
rect 451274 3340 451280 3392
rect 451332 3380 451338 3392
rect 452470 3380 452476 3392
rect 451332 3352 452476 3380
rect 451332 3340 451338 3352
rect 452470 3340 452476 3352
rect 452528 3340 452534 3392
rect 459554 3340 459560 3392
rect 459612 3380 459618 3392
rect 460842 3380 460848 3392
rect 459612 3352 460848 3380
rect 459612 3340 459618 3352
rect 460842 3340 460848 3352
rect 460900 3340 460906 3392
rect 502334 3340 502340 3392
rect 502392 3380 502398 3392
rect 503622 3380 503628 3392
rect 502392 3352 503628 3380
rect 502392 3340 502398 3352
rect 503622 3340 503628 3352
rect 503680 3340 503686 3392
rect 520274 3340 520280 3392
rect 520332 3380 520338 3392
rect 521470 3380 521476 3392
rect 520332 3352 521476 3380
rect 520332 3340 520338 3352
rect 521470 3340 521476 3352
rect 521528 3340 521534 3392
rect 536834 3340 536840 3392
rect 536892 3380 536898 3392
rect 538122 3380 538128 3392
rect 536892 3352 538128 3380
rect 536892 3340 536898 3352
rect 538122 3340 538128 3352
rect 538180 3340 538186 3392
rect 71866 3272 71872 3324
rect 71924 3312 71930 3324
rect 338574 3312 338580 3324
rect 71924 3284 338580 3312
rect 71924 3272 71930 3284
rect 338574 3272 338580 3284
rect 338632 3272 338638 3324
rect 64840 3216 71820 3244
rect 64840 3204 64846 3216
rect 76650 3204 76656 3256
rect 76708 3244 76714 3256
rect 77202 3244 77208 3256
rect 76708 3216 77208 3244
rect 76708 3204 76714 3216
rect 77202 3204 77208 3216
rect 77260 3204 77266 3256
rect 77846 3204 77852 3256
rect 77904 3244 77910 3256
rect 78582 3244 78588 3256
rect 77904 3216 78588 3244
rect 77904 3204 77910 3216
rect 78582 3204 78588 3216
rect 78640 3204 78646 3256
rect 80238 3204 80244 3256
rect 80296 3244 80302 3256
rect 81342 3244 81348 3256
rect 80296 3216 81348 3244
rect 80296 3204 80302 3216
rect 81342 3204 81348 3216
rect 81400 3204 81406 3256
rect 81434 3204 81440 3256
rect 81492 3244 81498 3256
rect 82538 3244 82544 3256
rect 81492 3216 82544 3244
rect 81492 3204 81498 3216
rect 82538 3204 82544 3216
rect 82596 3204 82602 3256
rect 339494 3244 339500 3256
rect 84856 3216 339500 3244
rect 55401 3179 55459 3185
rect 55401 3145 55413 3179
rect 55447 3176 55459 3179
rect 64509 3179 64567 3185
rect 64509 3176 64521 3179
rect 55447 3148 64521 3176
rect 55447 3145 55459 3148
rect 55401 3139 55459 3145
rect 64509 3145 64521 3148
rect 64555 3145 64567 3179
rect 64509 3139 64567 3145
rect 64877 3179 64935 3185
rect 64877 3145 64889 3179
rect 64923 3176 64935 3179
rect 74445 3179 74503 3185
rect 74445 3176 74457 3179
rect 64923 3148 74457 3176
rect 64923 3145 64935 3148
rect 64877 3139 64935 3145
rect 74445 3145 74457 3148
rect 74491 3145 74503 3179
rect 74445 3139 74503 3145
rect 79042 3136 79048 3188
rect 79100 3176 79106 3188
rect 84856 3176 84884 3216
rect 339494 3204 339500 3216
rect 339552 3204 339558 3256
rect 79100 3148 84884 3176
rect 79100 3136 79106 3148
rect 84930 3136 84936 3188
rect 84988 3176 84994 3188
rect 85482 3176 85488 3188
rect 84988 3148 85488 3176
rect 84988 3136 84994 3148
rect 85482 3136 85488 3148
rect 85540 3136 85546 3188
rect 86126 3136 86132 3188
rect 86184 3176 86190 3188
rect 86862 3176 86868 3188
rect 86184 3148 86868 3176
rect 86184 3136 86190 3148
rect 86862 3136 86868 3148
rect 86920 3136 86926 3188
rect 87322 3136 87328 3188
rect 87380 3176 87386 3188
rect 88242 3176 88248 3188
rect 87380 3148 88248 3176
rect 87380 3136 87386 3148
rect 88242 3136 88248 3148
rect 88300 3136 88306 3188
rect 88518 3136 88524 3188
rect 88576 3176 88582 3188
rect 89622 3176 89628 3188
rect 88576 3148 89628 3176
rect 88576 3136 88582 3148
rect 89622 3136 89628 3148
rect 89680 3136 89686 3188
rect 89714 3136 89720 3188
rect 89772 3176 89778 3188
rect 342714 3176 342720 3188
rect 89772 3148 342720 3176
rect 89772 3136 89778 3148
rect 342714 3136 342720 3148
rect 342772 3136 342778 3188
rect 344002 3108 344008 3120
rect 103900 3080 344008 3108
rect 20714 3000 20720 3052
rect 20772 3040 20778 3052
rect 22002 3040 22008 3052
rect 20772 3012 22008 3040
rect 20772 3000 20778 3012
rect 22002 3000 22008 3012
rect 22060 3000 22066 3052
rect 84197 3043 84255 3049
rect 84197 3009 84209 3043
rect 84243 3040 84255 3043
rect 84243 3012 93808 3040
rect 84243 3009 84255 3012
rect 84197 3003 84255 3009
rect 93780 2972 93808 3012
rect 96890 3000 96896 3052
rect 96948 3040 96954 3052
rect 103900 3040 103928 3080
rect 344002 3068 344008 3080
rect 344060 3068 344066 3120
rect 96948 3012 103928 3040
rect 96948 3000 96954 3012
rect 103974 3000 103980 3052
rect 104032 3040 104038 3052
rect 345382 3040 345388 3052
rect 104032 3012 345388 3040
rect 104032 3000 104038 3012
rect 345382 3000 345388 3012
rect 345440 3000 345446 3052
rect 99285 2975 99343 2981
rect 99285 2972 99297 2975
rect 93780 2944 99297 2972
rect 99285 2941 99297 2944
rect 99331 2941 99343 2975
rect 99285 2935 99343 2941
rect 119341 2975 119399 2981
rect 119341 2941 119353 2975
rect 119387 2972 119399 2975
rect 124125 2975 124183 2981
rect 124125 2972 124137 2975
rect 119387 2944 124137 2972
rect 119387 2941 119399 2944
rect 119341 2935 119399 2941
rect 124125 2941 124137 2944
rect 124171 2941 124183 2975
rect 124125 2935 124183 2941
rect 124217 2975 124275 2981
rect 124217 2941 124229 2975
rect 124263 2972 124275 2975
rect 348142 2972 348148 2984
rect 124263 2944 348148 2972
rect 124263 2941 124275 2944
rect 124217 2935 124275 2941
rect 348142 2932 348148 2944
rect 348200 2932 348206 2984
rect 34974 2864 34980 2916
rect 35032 2904 35038 2916
rect 35802 2904 35808 2916
rect 35032 2876 35808 2904
rect 35032 2864 35038 2876
rect 35802 2864 35808 2876
rect 35860 2864 35866 2916
rect 111150 2864 111156 2916
rect 111208 2904 111214 2916
rect 346670 2904 346676 2916
rect 111208 2876 346676 2904
rect 111208 2864 111214 2876
rect 346670 2864 346676 2876
rect 346728 2864 346734 2916
rect 92106 2796 92112 2848
rect 92164 2836 92170 2848
rect 92382 2836 92388 2848
rect 92164 2808 92388 2836
rect 92164 2796 92170 2808
rect 92382 2796 92388 2808
rect 92440 2796 92446 2848
rect 101493 2839 101551 2845
rect 101493 2805 101505 2839
rect 101539 2836 101551 2839
rect 117041 2839 117099 2845
rect 117041 2836 117053 2839
rect 101539 2808 117053 2836
rect 101539 2805 101551 2808
rect 101493 2799 101551 2805
rect 117041 2805 117053 2808
rect 117087 2805 117099 2839
rect 117041 2799 117099 2805
rect 117130 2796 117136 2848
rect 117188 2836 117194 2848
rect 347774 2836 347780 2848
rect 117188 2808 347780 2836
rect 117188 2796 117194 2808
rect 347774 2796 347780 2808
rect 347832 2796 347838 2848
rect 118234 2728 118240 2780
rect 118292 2768 118298 2780
rect 124217 2771 124275 2777
rect 124217 2768 124229 2771
rect 118292 2740 124229 2768
rect 118292 2728 118298 2740
rect 124217 2737 124229 2740
rect 124263 2737 124275 2771
rect 124217 2731 124275 2737
rect 267737 2771 267795 2777
rect 267737 2737 267749 2771
rect 267783 2768 267795 2771
rect 277305 2771 277363 2777
rect 277305 2768 277317 2771
rect 267783 2740 277317 2768
rect 267783 2737 267795 2740
rect 267737 2731 267795 2737
rect 277305 2737 277317 2740
rect 277351 2737 277363 2771
rect 277305 2731 277363 2737
rect 563054 2456 563060 2508
rect 563112 2496 563118 2508
rect 564342 2496 564348 2508
rect 563112 2468 564348 2496
rect 563112 2456 563118 2468
rect 564342 2456 564348 2468
rect 564400 2456 564406 2508
rect 356054 824 356060 876
rect 356112 864 356118 876
rect 357342 864 357348 876
rect 356112 836 357348 864
rect 356112 824 356118 836
rect 357342 824 357348 836
rect 357400 824 357406 876
rect 5258 552 5264 604
rect 5316 592 5322 604
rect 5442 592 5448 604
rect 5316 564 5448 592
rect 5316 552 5322 564
rect 5442 552 5448 564
rect 5500 552 5506 604
rect 90910 592 90916 604
rect 90871 564 90916 592
rect 90910 552 90916 564
rect 90968 552 90974 604
rect 100478 592 100484 604
rect 100439 564 100484 592
rect 100478 552 100484 564
rect 100536 552 100542 604
rect 107562 552 107568 604
rect 107620 592 107626 604
rect 107746 592 107752 604
rect 107620 564 107752 592
rect 107620 552 107626 564
rect 107746 552 107752 564
rect 107804 552 107810 604
rect 108758 592 108764 604
rect 108719 564 108764 592
rect 108758 552 108764 564
rect 108816 552 108822 604
rect 109954 552 109960 604
rect 110012 592 110018 604
rect 110322 592 110328 604
rect 110012 564 110328 592
rect 110012 552 110018 564
rect 110322 552 110328 564
rect 110380 552 110386 604
rect 280062 592 280068 604
rect 280023 564 280068 592
rect 280062 552 280068 564
rect 280120 552 280126 604
rect 324406 552 324412 604
rect 324464 592 324470 604
rect 325234 592 325240 604
rect 324464 564 325240 592
rect 324464 552 324470 564
rect 325234 552 325240 564
rect 325292 552 325298 604
rect 335354 552 335360 604
rect 335412 592 335418 604
rect 335906 592 335912 604
rect 335412 564 335912 592
rect 335412 552 335418 564
rect 335906 552 335912 564
rect 335964 552 335970 604
rect 336734 552 336740 604
rect 336792 592 336798 604
rect 337102 592 337108 604
rect 336792 564 337108 592
rect 336792 552 336798 564
rect 337102 552 337108 564
rect 337160 552 337166 604
rect 349154 552 349160 604
rect 349212 592 349218 604
rect 350258 592 350264 604
rect 349212 564 350264 592
rect 349212 552 349218 564
rect 350258 552 350264 564
rect 350316 552 350322 604
rect 394694 552 394700 604
rect 394752 592 394758 604
rect 395430 592 395436 604
rect 394752 564 395436 592
rect 394752 552 394758 564
rect 395430 552 395436 564
rect 395488 552 395494 604
rect 401594 552 401600 604
rect 401652 592 401658 604
rect 402514 592 402520 604
rect 401652 564 402520 592
rect 401652 552 401658 564
rect 402514 552 402520 564
rect 402572 552 402578 604
rect 402974 552 402980 604
rect 403032 592 403038 604
rect 403710 592 403716 604
rect 403032 564 403716 592
rect 403032 552 403038 564
rect 403710 552 403716 564
rect 403768 552 403774 604
rect 405734 552 405740 604
rect 405792 592 405798 604
rect 406102 592 406108 604
rect 405792 564 406108 592
rect 405792 552 405798 564
rect 406102 552 406108 564
rect 406160 552 406166 604
rect 409874 552 409880 604
rect 409932 592 409938 604
rect 410886 592 410892 604
rect 409932 564 410892 592
rect 409932 552 409938 564
rect 410886 552 410892 564
rect 410944 552 410950 604
rect 423674 552 423680 604
rect 423732 592 423738 604
rect 423950 592 423956 604
rect 423732 564 423956 592
rect 423732 552 423738 564
rect 423950 552 423956 564
rect 424008 552 424014 604
rect 426434 552 426440 604
rect 426492 592 426498 604
rect 427538 592 427544 604
rect 426492 564 427544 592
rect 426492 552 426498 564
rect 427538 552 427544 564
rect 427596 552 427602 604
rect 427814 552 427820 604
rect 427872 592 427878 604
rect 428734 592 428740 604
rect 427872 564 428740 592
rect 427872 552 427878 564
rect 428734 552 428740 564
rect 428792 552 428798 604
rect 430574 552 430580 604
rect 430632 592 430638 604
rect 431126 592 431132 604
rect 430632 564 431132 592
rect 430632 552 430638 564
rect 431126 552 431132 564
rect 431184 552 431190 604
rect 434714 552 434720 604
rect 434772 592 434778 604
rect 435818 592 435824 604
rect 434772 564 435824 592
rect 434772 552 434778 564
rect 435818 552 435824 564
rect 435876 552 435882 604
rect 436094 552 436100 604
rect 436152 592 436158 604
rect 437014 592 437020 604
rect 436152 564 437020 592
rect 436152 552 436158 564
rect 437014 552 437020 564
rect 437072 552 437078 604
rect 437474 552 437480 604
rect 437532 592 437538 604
rect 438210 592 438216 604
rect 437532 564 438216 592
rect 437532 552 437538 564
rect 438210 552 438216 564
rect 438268 552 438274 604
rect 438854 552 438860 604
rect 438912 592 438918 604
rect 439406 592 439412 604
rect 438912 564 439412 592
rect 438912 552 438918 564
rect 439406 552 439412 564
rect 439464 552 439470 604
rect 452654 552 452660 604
rect 452712 592 452718 604
rect 453666 592 453672 604
rect 452712 564 453672 592
rect 452712 552 452718 564
rect 453666 552 453672 564
rect 453724 552 453730 604
rect 455414 552 455420 604
rect 455472 592 455478 604
rect 456058 592 456064 604
rect 455472 564 456064 592
rect 455472 552 455478 564
rect 456058 552 456064 564
rect 456116 552 456122 604
rect 456794 552 456800 604
rect 456852 592 456858 604
rect 457254 592 457260 604
rect 456852 564 457260 592
rect 456852 552 456858 564
rect 457254 552 457260 564
rect 457312 552 457318 604
rect 462314 552 462320 604
rect 462372 592 462378 604
rect 463234 592 463240 604
rect 462372 564 463240 592
rect 462372 552 462378 564
rect 463234 552 463240 564
rect 463292 552 463298 604
rect 463694 552 463700 604
rect 463752 592 463758 604
rect 464430 592 464436 604
rect 463752 564 464436 592
rect 463752 552 463758 564
rect 464430 552 464436 564
rect 464488 552 464494 604
rect 466454 552 466460 604
rect 466512 592 466518 604
rect 466822 592 466828 604
rect 466512 564 466828 592
rect 466512 552 466518 564
rect 466822 552 466828 564
rect 466880 552 466886 604
rect 469214 552 469220 604
rect 469272 592 469278 604
rect 470318 592 470324 604
rect 469272 564 470324 592
rect 469272 552 469278 564
rect 470318 552 470324 564
rect 470376 552 470382 604
rect 470594 552 470600 604
rect 470652 592 470658 604
rect 471514 592 471520 604
rect 470652 564 471520 592
rect 470652 552 470658 564
rect 471514 552 471520 564
rect 471572 552 471578 604
rect 489914 552 489920 604
rect 489972 592 489978 604
rect 490558 592 490564 604
rect 489972 564 490564 592
rect 489972 552 489978 564
rect 490558 552 490564 564
rect 490616 552 490622 604
rect 495434 552 495440 604
rect 495492 592 495498 604
rect 496538 592 496544 604
rect 495492 564 496544 592
rect 495492 552 495498 564
rect 496538 552 496544 564
rect 496596 552 496602 604
rect 499574 552 499580 604
rect 499632 592 499638 604
rect 500126 592 500132 604
rect 499632 564 500132 592
rect 499632 552 499638 564
rect 500126 552 500132 564
rect 500184 552 500190 604
rect 506474 552 506480 604
rect 506532 592 506538 604
rect 507210 592 507216 604
rect 506532 564 507216 592
rect 506532 552 506538 564
rect 507210 552 507216 564
rect 507268 552 507274 604
rect 510614 552 510620 604
rect 510672 592 510678 604
rect 510798 592 510804 604
rect 510672 564 510804 592
rect 510672 552 510678 564
rect 510798 552 510804 564
rect 510856 552 510862 604
rect 513374 552 513380 604
rect 513432 592 513438 604
rect 514386 592 514392 604
rect 513432 564 514392 592
rect 513432 552 513438 564
rect 514386 552 514392 564
rect 514444 552 514450 604
rect 524414 552 524420 604
rect 524472 592 524478 604
rect 525058 592 525064 604
rect 524472 564 525064 592
rect 524472 552 524478 564
rect 525058 552 525064 564
rect 525116 552 525122 604
rect 538214 552 538220 604
rect 538272 592 538278 604
rect 539318 592 539324 604
rect 538272 564 539324 592
rect 538272 552 538278 564
rect 539318 552 539324 564
rect 539376 552 539382 604
rect 540974 552 540980 604
rect 541032 592 541038 604
rect 541710 592 541716 604
rect 541032 564 541716 592
rect 541032 552 541038 564
rect 541710 552 541716 564
rect 541768 552 541774 604
rect 542354 552 542360 604
rect 542412 592 542418 604
rect 542906 592 542912 604
rect 542412 564 542912 592
rect 542412 552 542418 564
rect 542906 552 542912 564
rect 542964 552 542970 604
rect 549254 552 549260 604
rect 549312 592 549318 604
rect 550082 592 550088 604
rect 549312 564 550088 592
rect 549312 552 549318 564
rect 550082 552 550088 564
rect 550140 552 550146 604
rect 556154 552 556160 604
rect 556212 592 556218 604
rect 557166 592 557172 604
rect 556212 564 557172 592
rect 556212 552 556218 564
rect 557166 552 557172 564
rect 557224 552 557230 604
<< via1 >>
rect 170312 700952 170364 701004
rect 293224 700952 293276 701004
rect 286968 700884 287020 700936
rect 413652 700884 413704 700936
rect 284208 700816 284260 700868
rect 429844 700816 429896 700868
rect 137836 700748 137888 700800
rect 294604 700748 294656 700800
rect 282828 700680 282880 700732
rect 462320 700680 462372 700732
rect 105452 700612 105504 700664
rect 295984 700612 296036 700664
rect 284116 700544 284168 700596
rect 478512 700544 478564 700596
rect 72976 700476 73028 700528
rect 297364 700476 297416 700528
rect 299480 700476 299532 700528
rect 300124 700476 300176 700528
rect 280068 700408 280120 700460
rect 527180 700408 527232 700460
rect 40500 700340 40552 700392
rect 300124 700340 300176 700392
rect 8116 700272 8168 700324
rect 301504 700272 301556 700324
rect 285588 700204 285640 700256
rect 397460 700204 397512 700256
rect 202788 700136 202840 700188
rect 291844 700136 291896 700188
rect 288348 700068 288400 700120
rect 364984 700068 365036 700120
rect 289728 700000 289780 700052
rect 348792 700000 348844 700052
rect 235172 699932 235224 699984
rect 290464 699932 290516 699984
rect 291108 699932 291160 699984
rect 299480 699932 299532 699984
rect 288256 699864 288308 699916
rect 332508 699864 332560 699916
rect 283840 699796 283892 699848
rect 291292 699796 291344 699848
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 89168 699660 89220 699712
rect 89628 699660 89680 699712
rect 542728 698232 542780 698284
rect 543556 698232 543608 698284
rect 275928 696940 275980 696992
rect 580172 696940 580224 696992
rect 154120 695512 154172 695564
rect 154212 695512 154264 695564
rect 218980 694152 219032 694204
rect 219164 694152 219216 694204
rect 219164 688644 219216 688696
rect 542728 688644 542780 688696
rect 154212 688576 154264 688628
rect 154396 688576 154448 688628
rect 219072 688576 219124 688628
rect 542544 688576 542596 688628
rect 559104 688576 559156 688628
rect 559656 688576 559708 688628
rect 277308 685856 277360 685908
rect 580172 685856 580224 685908
rect 154396 685788 154448 685840
rect 542452 684428 542504 684480
rect 559012 684428 559064 684480
rect 3516 681708 3568 681760
rect 305092 681708 305144 681760
rect 154304 676243 154356 676252
rect 154304 676209 154313 676243
rect 154313 676209 154347 676243
rect 154347 676209 154356 676243
rect 154304 676200 154356 676209
rect 218980 676175 219032 676184
rect 218980 676141 218989 676175
rect 218989 676141 219023 676175
rect 219023 676141 219032 676175
rect 218980 676132 219032 676141
rect 494060 676175 494112 676184
rect 494060 676141 494069 676175
rect 494069 676141 494103 676175
rect 494103 676141 494112 676175
rect 494060 676132 494112 676141
rect 154304 673480 154356 673532
rect 154488 673480 154540 673532
rect 274548 673480 274600 673532
rect 580172 673480 580224 673532
rect 3424 667904 3476 667956
rect 305644 667904 305696 667956
rect 219072 666544 219124 666596
rect 494152 666544 494204 666596
rect 542820 666544 542872 666596
rect 559380 666544 559432 666596
rect 219164 659608 219216 659660
rect 219348 659608 219400 659660
rect 219348 656820 219400 656872
rect 154304 654100 154356 654152
rect 154488 654100 154540 654152
rect 494060 654100 494112 654152
rect 494244 654100 494296 654152
rect 3056 652740 3108 652792
rect 306380 652740 306432 652792
rect 273168 650020 273220 650072
rect 580172 650020 580224 650072
rect 219256 647275 219308 647284
rect 219256 647241 219265 647275
rect 219265 647241 219299 647275
rect 219299 647241 219308 647275
rect 219256 647232 219308 647241
rect 542544 647232 542596 647284
rect 542636 647232 542688 647284
rect 559104 647232 559156 647284
rect 559196 647232 559248 647284
rect 219256 640364 219308 640416
rect 542544 640364 542596 640416
rect 542636 640364 542688 640416
rect 559104 640364 559156 640416
rect 559196 640364 559248 640416
rect 219072 640228 219124 640280
rect 274456 638936 274508 638988
rect 580172 638936 580224 638988
rect 219072 637508 219124 637560
rect 219164 637508 219216 637560
rect 154304 634788 154356 634840
rect 154488 634788 154540 634840
rect 494060 634788 494112 634840
rect 494244 634788 494296 634840
rect 542452 630640 542504 630692
rect 542636 630640 542688 630692
rect 559012 630640 559064 630692
rect 559196 630640 559248 630692
rect 271788 626560 271840 626612
rect 580172 626560 580224 626612
rect 219348 626535 219400 626544
rect 219348 626501 219357 626535
rect 219357 626501 219391 626535
rect 219391 626501 219400 626535
rect 219348 626492 219400 626501
rect 3424 623772 3476 623824
rect 309140 623772 309192 623824
rect 219348 616879 219400 616888
rect 219348 616845 219357 616879
rect 219357 616845 219391 616879
rect 219391 616845 219400 616879
rect 219348 616836 219400 616845
rect 154304 615476 154356 615528
rect 154488 615476 154540 615528
rect 494060 615476 494112 615528
rect 494244 615476 494296 615528
rect 219348 611396 219400 611448
rect 542452 611328 542504 611380
rect 542636 611328 542688 611380
rect 559012 611328 559064 611380
rect 559196 611328 559248 611380
rect 3424 609968 3476 610020
rect 308404 609968 308456 610020
rect 219072 608719 219124 608728
rect 219072 608685 219081 608719
rect 219081 608685 219115 608719
rect 219115 608685 219124 608719
rect 219072 608676 219124 608685
rect 219072 608540 219124 608592
rect 542544 608583 542596 608592
rect 542544 608549 542553 608583
rect 542553 608549 542587 608583
rect 542587 608549 542596 608583
rect 542544 608540 542596 608549
rect 559104 608583 559156 608592
rect 559104 608549 559113 608583
rect 559113 608549 559147 608583
rect 559147 608549 559156 608583
rect 559104 608540 559156 608549
rect 270408 603100 270460 603152
rect 580172 603100 580224 603152
rect 542728 601672 542780 601724
rect 559288 601672 559340 601724
rect 219256 601579 219308 601588
rect 219256 601545 219265 601579
rect 219265 601545 219299 601579
rect 219299 601545 219308 601579
rect 219256 601536 219308 601545
rect 219256 598884 219308 598936
rect 542728 598927 542780 598936
rect 542728 598893 542737 598927
rect 542737 598893 542771 598927
rect 542771 598893 542780 598927
rect 542728 598884 542780 598893
rect 559288 598927 559340 598936
rect 559288 598893 559297 598927
rect 559297 598893 559331 598927
rect 559331 598893 559340 598927
rect 559288 598884 559340 598893
rect 154304 596164 154356 596216
rect 154488 596164 154540 596216
rect 494060 596164 494112 596216
rect 494244 596164 494296 596216
rect 3240 594804 3292 594856
rect 309232 594804 309284 594856
rect 270316 592016 270368 592068
rect 580172 592016 580224 592068
rect 219164 589339 219216 589348
rect 219164 589305 219173 589339
rect 219173 589305 219207 589339
rect 219207 589305 219216 589339
rect 219164 589296 219216 589305
rect 542820 589296 542872 589348
rect 559380 589296 559432 589348
rect 154304 589271 154356 589280
rect 154304 589237 154313 589271
rect 154313 589237 154347 589271
rect 154347 589237 154356 589271
rect 154304 589228 154356 589237
rect 493876 589228 493928 589280
rect 494152 589228 494204 589280
rect 218980 582360 219032 582412
rect 219164 582360 219216 582412
rect 542820 582428 542872 582480
rect 559380 582428 559432 582480
rect 542728 582292 542780 582344
rect 559288 582292 559340 582344
rect 154304 579751 154356 579760
rect 154304 579717 154313 579751
rect 154313 579717 154347 579751
rect 154347 579717 154356 579751
rect 154304 579708 154356 579717
rect 269028 579640 269080 579692
rect 580172 579640 580224 579692
rect 154212 579572 154264 579624
rect 154396 579572 154448 579624
rect 218980 579572 219032 579624
rect 218888 569959 218940 569968
rect 218888 569925 218897 569959
rect 218897 569925 218931 569959
rect 218931 569925 218940 569959
rect 218888 569916 218940 569925
rect 494152 569891 494204 569900
rect 494152 569857 494161 569891
rect 494161 569857 494195 569891
rect 494195 569857 494204 569891
rect 494152 569848 494204 569857
rect 3424 567196 3476 567248
rect 311900 567196 311952 567248
rect 542452 563116 542504 563168
rect 559012 563116 559064 563168
rect 218888 563048 218940 563100
rect 494336 563048 494388 563100
rect 154212 562912 154264 562964
rect 154396 562912 154448 562964
rect 542452 562980 542504 563032
rect 559012 562980 559064 563032
rect 218980 562912 219032 562964
rect 542452 560235 542504 560244
rect 542452 560201 542461 560235
rect 542461 560201 542495 560235
rect 542495 560201 542504 560235
rect 542452 560192 542504 560201
rect 559012 560235 559064 560244
rect 559012 560201 559021 560235
rect 559021 560201 559055 560235
rect 559055 560201 559064 560235
rect 559012 560192 559064 560201
rect 266268 556180 266320 556232
rect 580172 556180 580224 556232
rect 218888 553435 218940 553444
rect 218888 553401 218897 553435
rect 218897 553401 218931 553435
rect 218931 553401 218940 553435
rect 218888 553392 218940 553401
rect 3148 552032 3200 552084
rect 311164 552032 311216 552084
rect 218888 550647 218940 550656
rect 218888 550613 218897 550647
rect 218897 550613 218931 550647
rect 218931 550613 218940 550647
rect 218888 550604 218940 550613
rect 494152 550604 494204 550656
rect 494428 550604 494480 550656
rect 542636 550604 542688 550656
rect 559196 550604 559248 550656
rect 267556 545096 267608 545148
rect 580172 545096 580224 545148
rect 218888 543736 218940 543788
rect 494428 543804 494480 543856
rect 494336 543668 494388 543720
rect 218980 543600 219032 543652
rect 542452 543600 542504 543652
rect 542636 543600 542688 543652
rect 559012 543600 559064 543652
rect 559196 543600 559248 543652
rect 3424 538228 3476 538280
rect 313372 538228 313424 538280
rect 542452 534012 542504 534064
rect 542636 534012 542688 534064
rect 559012 534012 559064 534064
rect 559196 534012 559248 534064
rect 266176 532720 266228 532772
rect 580172 532720 580224 532772
rect 494152 531292 494204 531344
rect 494428 531292 494480 531344
rect 154396 531267 154448 531276
rect 154396 531233 154405 531267
rect 154405 531233 154439 531267
rect 154439 531233 154448 531267
rect 154396 531224 154448 531233
rect 494428 524492 494480 524544
rect 542636 524424 542688 524476
rect 559196 524424 559248 524476
rect 494336 524356 494388 524408
rect 542728 524356 542780 524408
rect 559288 524356 559340 524408
rect 218980 524288 219032 524340
rect 219164 524288 219216 524340
rect 154488 521636 154540 521688
rect 218796 514632 218848 514684
rect 219072 514632 219124 514684
rect 494152 511980 494204 512032
rect 494428 511980 494480 512032
rect 542544 511980 542596 512032
rect 542820 511980 542872 512032
rect 559104 511980 559156 512032
rect 559380 511980 559432 512032
rect 154396 511955 154448 511964
rect 154396 511921 154405 511955
rect 154405 511921 154439 511955
rect 154439 511921 154448 511955
rect 154396 511912 154448 511921
rect 219072 510595 219124 510604
rect 219072 510561 219081 510595
rect 219081 510561 219115 510595
rect 219115 510561 219124 510595
rect 219072 510552 219124 510561
rect 3424 509328 3476 509380
rect 314660 509328 314712 509380
rect 263508 509260 263560 509312
rect 580172 509260 580224 509312
rect 219072 505087 219124 505096
rect 219072 505053 219081 505087
rect 219081 505053 219115 505087
rect 219115 505053 219124 505087
rect 219072 505044 219124 505053
rect 154488 502324 154540 502376
rect 494244 502324 494296 502376
rect 494428 502324 494480 502376
rect 542636 502324 542688 502376
rect 542820 502324 542872 502376
rect 559196 502324 559248 502376
rect 559380 502324 559432 502376
rect 264888 498176 264940 498228
rect 580172 498176 580224 498228
rect 3424 495456 3476 495508
rect 313924 495456 313976 495508
rect 219072 492668 219124 492720
rect 219164 492668 219216 492720
rect 542544 492643 542596 492652
rect 542544 492609 542553 492643
rect 542553 492609 542587 492643
rect 542587 492609 542596 492643
rect 542544 492600 542596 492609
rect 559104 492643 559156 492652
rect 559104 492609 559113 492643
rect 559113 492609 559147 492643
rect 559147 492609 559156 492643
rect 559104 492600 559156 492609
rect 154304 485800 154356 485852
rect 219164 485800 219216 485852
rect 262128 485800 262180 485852
rect 580172 485800 580224 485852
rect 154396 485664 154448 485716
rect 542544 485775 542596 485784
rect 542544 485741 542553 485775
rect 542553 485741 542587 485775
rect 542587 485741 542596 485775
rect 542544 485732 542596 485741
rect 559104 485775 559156 485784
rect 559104 485741 559113 485775
rect 559113 485741 559147 485775
rect 559147 485741 559156 485775
rect 559104 485732 559156 485741
rect 219256 485664 219308 485716
rect 154396 482987 154448 482996
rect 154396 482953 154405 482987
rect 154405 482953 154439 482987
rect 154439 482953 154448 482987
rect 154396 482944 154448 482953
rect 3148 480224 3200 480276
rect 316040 480224 316092 480276
rect 494060 480224 494112 480276
rect 494244 480224 494296 480276
rect 219072 476076 219124 476128
rect 219256 476076 219308 476128
rect 542452 476076 542504 476128
rect 542636 476076 542688 476128
rect 559012 476076 559064 476128
rect 559196 476076 559248 476128
rect 154396 476051 154448 476060
rect 154396 476017 154405 476051
rect 154405 476017 154439 476051
rect 154439 476017 154448 476051
rect 154396 476008 154448 476017
rect 542636 466488 542688 466540
rect 559196 466488 559248 466540
rect 542544 463743 542596 463752
rect 542544 463709 542553 463743
rect 542553 463709 542587 463743
rect 542587 463709 542596 463743
rect 542544 463700 542596 463709
rect 559104 463743 559156 463752
rect 559104 463709 559113 463743
rect 559113 463709 559147 463743
rect 559147 463709 559156 463743
rect 559104 463700 559156 463709
rect 291384 463632 291436 463684
rect 291844 463632 291896 463684
rect 294512 463632 294564 463684
rect 297364 463632 297416 463684
rect 300860 463632 300912 463684
rect 301504 463632 301556 463684
rect 303988 463632 304040 463684
rect 308404 463632 308456 463684
rect 311348 463632 311400 463684
rect 290464 463564 290516 463616
rect 293500 463564 293552 463616
rect 298744 463564 298796 463616
rect 300124 463564 300176 463616
rect 302976 463564 303028 463616
rect 311164 463564 311216 463616
rect 314568 463564 314620 463616
rect 280896 463496 280948 463548
rect 267648 463428 267700 463480
rect 295616 463428 295668 463480
rect 295984 463428 296036 463480
rect 299756 463428 299808 463480
rect 219072 463360 219124 463412
rect 293224 463360 293276 463412
rect 296628 463360 296680 463412
rect 129740 463292 129792 463344
rect 154304 463292 154356 463344
rect 294604 463292 294656 463344
rect 297732 463292 297784 463344
rect 129832 463224 129884 463276
rect 89628 463088 89680 463140
rect 147680 463156 147732 463208
rect 301872 463224 301924 463276
rect 147772 463088 147824 463140
rect 279792 463156 279844 463208
rect 277676 463088 277728 463140
rect 281908 463156 281960 463208
rect 282828 463156 282880 463208
rect 282920 463156 282972 463208
rect 284116 463156 284168 463208
rect 286140 463156 286192 463208
rect 286968 463156 287020 463208
rect 287152 463156 287204 463208
rect 288348 463156 288400 463208
rect 290372 463156 290424 463208
rect 291108 463156 291160 463208
rect 494244 463156 494296 463208
rect 24768 463020 24820 463072
rect 264060 462952 264112 463004
rect 264888 462952 264940 463004
rect 265072 462952 265124 463004
rect 266176 462952 266228 463004
rect 268200 462952 268252 463004
rect 269028 462952 269080 463004
rect 269304 462952 269356 463004
rect 270408 462952 270460 463004
rect 272432 462952 272484 463004
rect 273168 462952 273220 463004
rect 273444 462952 273496 463004
rect 274456 462952 274508 463004
rect 278780 462952 278832 463004
rect 280068 462952 280120 463004
rect 542544 463088 542596 463140
rect 305000 463020 305052 463072
rect 305644 463020 305696 463072
rect 308220 463020 308272 463072
rect 313924 463020 313976 463072
rect 317696 463020 317748 463072
rect 559104 462952 559156 463004
rect 31024 462884 31076 462936
rect 342904 462884 342956 462936
rect 4620 462816 4672 462868
rect 320824 462816 320876 462868
rect 2964 462748 3016 462800
rect 319812 462748 319864 462800
rect 3240 462680 3292 462732
rect 322940 462680 322992 462732
rect 3148 462612 3200 462664
rect 324044 462612 324096 462664
rect 259828 462544 259880 462596
rect 580080 462544 580132 462596
rect 238760 462476 238812 462528
rect 577504 462476 577556 462528
rect 236644 462408 236696 462460
rect 580356 462408 580408 462460
rect 3424 462340 3476 462392
rect 348240 462340 348292 462392
rect 260840 460232 260892 460284
rect 580172 460232 580224 460284
rect 4712 460164 4764 460216
rect 327172 460164 327224 460216
rect 5448 460096 5500 460148
rect 330300 460096 330352 460148
rect 5264 460028 5316 460080
rect 333060 460028 333112 460080
rect 250720 459960 250772 460012
rect 579988 459960 580040 460012
rect 5080 459892 5132 459944
rect 336372 459892 336424 459944
rect 247592 459824 247644 459876
rect 579712 459824 579764 459876
rect 4896 459756 4948 459808
rect 339500 459756 339552 459808
rect 244096 459688 244148 459740
rect 580816 459688 580868 459740
rect 241152 459620 241204 459672
rect 580632 459620 580684 459672
rect 235908 459552 235960 459604
rect 580264 459552 580316 459604
rect 238024 459459 238076 459468
rect 238024 459425 238033 459459
rect 238033 459425 238067 459459
rect 238067 459425 238076 459459
rect 238024 459416 238076 459425
rect 240048 459459 240100 459468
rect 240048 459425 240057 459459
rect 240057 459425 240091 459459
rect 240091 459425 240100 459459
rect 240048 459416 240100 459425
rect 243360 459459 243412 459468
rect 243360 459425 243369 459459
rect 243369 459425 243403 459459
rect 243403 459425 243412 459459
rect 243360 459416 243412 459425
rect 246488 459459 246540 459468
rect 246488 459425 246497 459459
rect 246497 459425 246531 459459
rect 246531 459425 246540 459459
rect 246488 459416 246540 459425
rect 249616 459459 249668 459468
rect 249616 459425 249625 459459
rect 249625 459425 249659 459459
rect 249659 459425 249668 459459
rect 249616 459416 249668 459425
rect 254952 459459 255004 459468
rect 254952 459425 254961 459459
rect 254961 459425 254995 459459
rect 254995 459425 255004 459459
rect 254952 459416 255004 459425
rect 257988 459416 258040 459468
rect 349896 459416 349948 459468
rect 3056 459348 3108 459400
rect 321652 459348 321704 459400
rect 4068 459280 4120 459332
rect 325884 459280 325936 459332
rect 329012 459348 329064 459400
rect 327908 459280 327960 459332
rect 331220 459323 331272 459332
rect 331220 459289 331229 459323
rect 331229 459289 331263 459323
rect 331263 459289 331272 459323
rect 331220 459280 331272 459289
rect 332140 459323 332192 459332
rect 332140 459289 332149 459323
rect 332149 459289 332183 459323
rect 332183 459289 332192 459323
rect 332140 459280 332192 459289
rect 334164 459323 334216 459332
rect 334164 459289 334173 459323
rect 334173 459289 334207 459323
rect 334207 459289 334216 459323
rect 334164 459280 334216 459289
rect 335360 459323 335412 459332
rect 335360 459289 335369 459323
rect 335369 459289 335403 459323
rect 335403 459289 335412 459323
rect 337292 459323 337344 459332
rect 335360 459280 335412 459289
rect 337292 459289 337301 459323
rect 337301 459289 337335 459323
rect 337335 459289 337344 459323
rect 337292 459280 337344 459289
rect 338396 459323 338448 459332
rect 338396 459289 338405 459323
rect 338405 459289 338439 459323
rect 338439 459289 338448 459323
rect 338396 459280 338448 459289
rect 340696 459323 340748 459332
rect 340696 459289 340705 459323
rect 340705 459289 340739 459323
rect 340739 459289 340748 459323
rect 340696 459280 340748 459289
rect 341524 459323 341576 459332
rect 341524 459289 341533 459323
rect 341533 459289 341567 459323
rect 341567 459289 341576 459323
rect 341524 459280 341576 459289
rect 3976 459144 4028 459196
rect 5356 459076 5408 459128
rect 579896 459076 579948 459128
rect 5172 459008 5224 459060
rect 3884 458940 3936 458992
rect 3792 458872 3844 458924
rect 580080 458804 580132 458856
rect 4988 458736 5040 458788
rect 3700 458668 3752 458720
rect 4804 458600 4856 458652
rect 580908 458532 580960 458584
rect 580724 458464 580776 458516
rect 3608 458396 3660 458448
rect 3516 458328 3568 458380
rect 580540 458260 580592 458312
rect 580448 458192 580500 458244
rect 579712 451596 579764 451648
rect 580172 451596 580224 451648
rect 2780 437996 2832 438048
rect 4620 437996 4672 438048
rect 349896 405628 349948 405680
rect 579804 405628 579856 405680
rect 281724 340144 281776 340196
rect 282460 340144 282512 340196
rect 299572 340144 299624 340196
rect 300584 340144 300636 340196
rect 317972 340144 318024 340196
rect 262588 339056 262640 339108
rect 263048 339056 263100 339108
rect 270684 339056 270736 339108
rect 271144 339056 271196 339108
rect 302976 339056 303028 339108
rect 303344 339056 303396 339108
rect 243360 338920 243412 338972
rect 243728 338920 243780 338972
rect 267740 338920 267792 338972
rect 268200 338920 268252 338972
rect 309140 338920 309192 338972
rect 309508 338920 309560 338972
rect 316500 338920 316552 338972
rect 316868 338920 316920 338972
rect 258724 338852 258776 338904
rect 259092 338852 259144 338904
rect 232872 338784 232924 338836
rect 233148 338784 233200 338836
rect 241704 338784 241756 338836
rect 242072 338784 242124 338836
rect 231860 338648 231912 338700
rect 232136 338648 232188 338700
rect 238024 338648 238076 338700
rect 238300 338648 238352 338700
rect 259460 338648 259512 338700
rect 259828 338648 259880 338700
rect 343732 338648 343784 338700
rect 344100 338648 344152 338700
rect 242992 338512 243044 338564
rect 243268 338512 243320 338564
rect 334164 338512 334216 338564
rect 334532 338512 334584 338564
rect 272156 338376 272208 338428
rect 272616 338376 272668 338428
rect 280252 338376 280304 338428
rect 280620 338376 280672 338428
rect 287244 338376 287296 338428
rect 287704 338376 287756 338428
rect 290004 338376 290056 338428
rect 290280 338376 290332 338428
rect 341064 338376 341116 338428
rect 341340 338376 341392 338428
rect 309876 338104 309928 338156
rect 310060 338104 310112 338156
rect 317880 338147 317932 338156
rect 317880 338113 317889 338147
rect 317889 338113 317923 338147
rect 317923 338113 317932 338147
rect 317880 338104 317932 338113
rect 319536 338104 319588 338156
rect 320088 338104 320140 338156
rect 86868 338036 86920 338088
rect 341616 338036 341668 338088
rect 93768 337968 93820 338020
rect 343088 337968 343140 338020
rect 82728 337900 82780 337952
rect 340880 337900 340932 337952
rect 75828 337832 75880 337884
rect 339408 337832 339460 337884
rect 62028 337764 62080 337816
rect 336464 337764 336516 337816
rect 68928 337696 68980 337748
rect 337936 337696 337988 337748
rect 57888 337628 57940 337680
rect 335728 337628 335780 337680
rect 44088 337560 44140 337612
rect 55128 337492 55180 337544
rect 42708 337424 42760 337476
rect 35808 337356 35860 337408
rect 322020 337356 322072 337408
rect 322204 337356 322256 337408
rect 322756 337356 322808 337408
rect 323124 337424 323176 337476
rect 323768 337424 323820 337476
rect 323952 337424 324004 337476
rect 330944 337492 330996 337544
rect 332784 337492 332836 337544
rect 334992 337424 335044 337476
rect 332600 337356 332652 337408
rect 100668 337288 100720 337340
rect 344560 337288 344612 337340
rect 107476 337220 107528 337272
rect 346032 337220 346084 337272
rect 115848 337152 115900 337204
rect 347504 337152 347556 337204
rect 122748 337084 122800 337136
rect 348976 337084 349028 337136
rect 173164 337016 173216 337068
rect 345756 337016 345808 337068
rect 182824 336948 182876 337000
rect 347228 336948 347280 337000
rect 186964 336880 187016 336932
rect 348700 336880 348752 336932
rect 191104 336812 191156 336864
rect 349436 336812 349488 336864
rect 195244 336744 195296 336796
rect 349712 336744 349764 336796
rect 107476 336719 107528 336728
rect 107476 336685 107485 336719
rect 107485 336685 107519 336719
rect 107519 336685 107528 336719
rect 107476 336676 107528 336685
rect 271972 336676 272024 336728
rect 272156 336676 272208 336728
rect 279516 336719 279568 336728
rect 279516 336685 279525 336719
rect 279525 336685 279559 336719
rect 279559 336685 279568 336719
rect 279516 336676 279568 336685
rect 305368 336676 305420 336728
rect 305552 336676 305604 336728
rect 291384 336608 291436 336660
rect 291752 336608 291804 336660
rect 313372 335996 313424 336048
rect 313648 335996 313700 336048
rect 313556 335928 313608 335980
rect 320180 335928 320232 335980
rect 320824 335928 320876 335980
rect 236000 335860 236052 335912
rect 236460 335860 236512 335912
rect 236184 335792 236236 335844
rect 236644 335792 236696 335844
rect 245752 335792 245804 335844
rect 245936 335792 245988 335844
rect 261300 335792 261352 335844
rect 269212 335792 269264 335844
rect 270224 335792 270276 335844
rect 273444 335792 273496 335844
rect 273628 335792 273680 335844
rect 299664 335792 299716 335844
rect 299848 335792 299900 335844
rect 311992 335792 312044 335844
rect 312544 335792 312596 335844
rect 232228 335724 232280 335776
rect 317696 335792 317748 335844
rect 317972 335792 318024 335844
rect 284484 335724 284536 335776
rect 284668 335724 284720 335776
rect 291292 335724 291344 335776
rect 292304 335724 292356 335776
rect 303804 335724 303856 335776
rect 303988 335724 304040 335776
rect 313556 335724 313608 335776
rect 328552 335724 328604 335776
rect 328828 335724 328880 335776
rect 233332 335656 233384 335708
rect 234252 335656 234304 335708
rect 237380 335656 237432 335708
rect 238392 335656 238444 335708
rect 247040 335656 247092 335708
rect 248144 335656 248196 335708
rect 248420 335656 248472 335708
rect 248880 335656 248932 335708
rect 249892 335656 249944 335708
rect 250352 335656 250404 335708
rect 251364 335656 251416 335708
rect 251824 335656 251876 335708
rect 252652 335656 252704 335708
rect 253296 335656 253348 335708
rect 254308 335656 254360 335708
rect 254492 335656 254544 335708
rect 255504 335656 255556 335708
rect 256056 335656 256108 335708
rect 261300 335656 261352 335708
rect 262220 335656 262272 335708
rect 263324 335656 263376 335708
rect 266636 335656 266688 335708
rect 267556 335656 267608 335708
rect 267832 335656 267884 335708
rect 268752 335656 268804 335708
rect 269304 335656 269356 335708
rect 270224 335656 270276 335708
rect 276204 335656 276256 335708
rect 277308 335656 277360 335708
rect 277400 335656 277452 335708
rect 278228 335656 278280 335708
rect 280160 335656 280212 335708
rect 281264 335656 281316 335708
rect 281540 335656 281592 335708
rect 282736 335656 282788 335708
rect 284392 335656 284444 335708
rect 284944 335656 284996 335708
rect 286048 335656 286100 335708
rect 286784 335656 286836 335708
rect 289912 335656 289964 335708
rect 290740 335656 290792 335708
rect 291568 335656 291620 335708
rect 292028 335656 292080 335708
rect 293040 335656 293092 335708
rect 293684 335656 293736 335708
rect 296812 335656 296864 335708
rect 297456 335656 297508 335708
rect 307760 335656 307812 335708
rect 308588 335656 308640 335708
rect 310980 335656 311032 335708
rect 311716 335656 311768 335708
rect 313648 335656 313700 335708
rect 314200 335656 314252 335708
rect 314752 335656 314804 335708
rect 315856 335656 315908 335708
rect 324320 335656 324372 335708
rect 325056 335656 325108 335708
rect 325792 335656 325844 335708
rect 326252 335656 326304 335708
rect 328460 335656 328512 335708
rect 329012 335656 329064 335708
rect 338304 335656 338356 335708
rect 338764 335656 338816 335708
rect 339500 335656 339552 335708
rect 339960 335656 340012 335708
rect 342720 335656 342772 335708
rect 342904 335656 342956 335708
rect 345204 335656 345256 335708
rect 346124 335656 346176 335708
rect 348056 335656 348108 335708
rect 348332 335656 348384 335708
rect 229192 335588 229244 335640
rect 230112 335588 230164 335640
rect 231952 335588 232004 335640
rect 232228 335588 232280 335640
rect 233240 335588 233292 335640
rect 233516 335588 233568 335640
rect 234712 335588 234764 335640
rect 234988 335588 235040 335640
rect 235172 335588 235224 335640
rect 235724 335588 235776 335640
rect 237472 335588 237524 335640
rect 237932 335588 237984 335640
rect 239128 335588 239180 335640
rect 239864 335588 239916 335640
rect 240416 335588 240468 335640
rect 241060 335588 241112 335640
rect 241612 335588 241664 335640
rect 242348 335588 242400 335640
rect 244280 335588 244332 335640
rect 245200 335588 245252 335640
rect 247500 335588 247552 335640
rect 247960 335588 248012 335640
rect 248696 335588 248748 335640
rect 249432 335588 249484 335640
rect 250168 335588 250220 335640
rect 250904 335588 250956 335640
rect 251640 335588 251692 335640
rect 252100 335588 252152 335640
rect 252560 335588 252612 335640
rect 253112 335588 253164 335640
rect 254124 335588 254176 335640
rect 254768 335588 254820 335640
rect 255780 335588 255832 335640
rect 256240 335588 256292 335640
rect 257344 335588 257396 335640
rect 257712 335588 257764 335640
rect 258632 335588 258684 335640
rect 259184 335588 259236 335640
rect 259644 335588 259696 335640
rect 260380 335588 260432 335640
rect 261208 335588 261260 335640
rect 261668 335588 261720 335640
rect 262404 335588 262456 335640
rect 262680 335588 262732 335640
rect 263968 335588 264020 335640
rect 264888 335588 264940 335640
rect 265164 335588 265216 335640
rect 265348 335588 265400 335640
rect 266360 335588 266412 335640
rect 266820 335588 266872 335640
rect 268384 335588 268436 335640
rect 269028 335588 269080 335640
rect 269672 335588 269724 335640
rect 270408 335588 270460 335640
rect 270500 335588 270552 335640
rect 271604 335588 271656 335640
rect 272064 335588 272116 335640
rect 273168 335588 273220 335640
rect 273720 335588 273772 335640
rect 274548 335588 274600 335640
rect 276112 335588 276164 335640
rect 276572 335588 276624 335640
rect 277768 335588 277820 335640
rect 278320 335588 278372 335640
rect 280344 335588 280396 335640
rect 280712 335588 280764 335640
rect 282276 335588 282328 335640
rect 282828 335588 282880 335640
rect 283288 335588 283340 335640
rect 283932 335588 283984 335640
rect 285680 335588 285732 335640
rect 286416 335588 286468 335640
rect 287612 335588 287664 335640
rect 288072 335588 288124 335640
rect 288532 335588 288584 335640
rect 289084 335588 289136 335640
rect 289820 335588 289872 335640
rect 290556 335588 290608 335640
rect 291476 335588 291528 335640
rect 291844 335588 291896 335640
rect 292948 335588 293000 335640
rect 293500 335588 293552 335640
rect 298468 335588 298520 335640
rect 299112 335588 299164 335640
rect 302608 335588 302660 335640
rect 303436 335588 303488 335640
rect 303988 335588 304040 335640
rect 304540 335588 304592 335640
rect 305184 335588 305236 335640
rect 305736 335588 305788 335640
rect 306656 335588 306708 335640
rect 306932 335588 306984 335640
rect 307944 335588 307996 335640
rect 308680 335588 308732 335640
rect 310520 335588 310572 335640
rect 310704 335588 310756 335640
rect 312176 335588 312228 335640
rect 313188 335588 313240 335640
rect 313280 335588 313332 335640
rect 314292 335588 314344 335640
rect 316132 335588 316184 335640
rect 316960 335588 317012 335640
rect 318984 335588 319036 335640
rect 319444 335588 319496 335640
rect 320640 335588 320692 335640
rect 321100 335588 321152 335640
rect 324780 335588 324832 335640
rect 325332 335588 325384 335640
rect 325884 335588 325936 335640
rect 326344 335588 326396 335640
rect 327264 335588 327316 335640
rect 327540 335588 327592 335640
rect 329932 335588 329984 335640
rect 330484 335588 330536 335640
rect 331404 335588 331456 335640
rect 332140 335588 332192 335640
rect 332692 335588 332744 335640
rect 333428 335588 333480 335640
rect 334348 335588 334400 335640
rect 334624 335588 334676 335640
rect 337016 335588 337068 335640
rect 337568 335588 337620 335640
rect 338488 335588 338540 335640
rect 339040 335588 339092 335640
rect 339776 335588 339828 335640
rect 340512 335588 340564 335640
rect 340972 335588 341024 335640
rect 341708 335588 341760 335640
rect 342444 335588 342496 335640
rect 343180 335588 343232 335640
rect 343916 335588 343968 335640
rect 344192 335588 344244 335640
rect 345020 335588 345072 335640
rect 345664 335588 345716 335640
rect 347780 335588 347832 335640
rect 348424 335588 348476 335640
rect 248512 335520 248564 335572
rect 249156 335520 249208 335572
rect 249984 335520 250036 335572
rect 250628 335520 250680 335572
rect 251456 335520 251508 335572
rect 252376 335520 252428 335572
rect 277584 335520 277636 335572
rect 278504 335520 278556 335572
rect 287152 335520 287204 335572
rect 287980 335520 288032 335572
rect 291292 335520 291344 335572
rect 292212 335520 292264 335572
rect 292764 335520 292816 335572
rect 293408 335520 293460 335572
rect 312084 335520 312136 335572
rect 312636 335520 312688 335572
rect 317788 335520 317840 335572
rect 318064 335520 318116 335572
rect 345112 335520 345164 335572
rect 345388 335520 345440 335572
rect 233516 335452 233568 335504
rect 233976 335452 234028 335504
rect 234988 335452 235040 335504
rect 235448 335452 235500 335504
rect 243084 335452 243136 335504
rect 244004 335452 244056 335504
rect 258172 335452 258224 335504
rect 259000 335452 259052 335504
rect 262404 335452 262456 335504
rect 263140 335452 263192 335504
rect 266820 335452 266872 335504
rect 267372 335452 267424 335504
rect 276112 335452 276164 335504
rect 276664 335452 276716 335504
rect 311072 335452 311124 335504
rect 311624 335452 311676 335504
rect 315028 335452 315080 335504
rect 315304 335452 315356 335504
rect 327356 335452 327408 335504
rect 327540 335452 327592 335504
rect 342536 335452 342588 335504
rect 343456 335452 343508 335504
rect 238852 335384 238904 335436
rect 239220 335384 239272 335436
rect 258632 335384 258684 335436
rect 259276 335384 259328 335436
rect 320916 335384 320968 335436
rect 321468 335384 321520 335436
rect 296996 335316 297048 335368
rect 297916 335316 297968 335368
rect 327356 335316 327408 335368
rect 328276 335316 328328 335368
rect 238852 335248 238904 335300
rect 239588 335248 239640 335300
rect 269764 335180 269816 335232
rect 270132 335180 270184 335232
rect 320180 335180 320232 335232
rect 325884 335180 325936 335232
rect 326528 335180 326580 335232
rect 265072 334976 265124 335028
rect 266176 334976 266228 335028
rect 323308 334976 323360 335028
rect 324044 334976 324096 335028
rect 275652 334704 275704 334756
rect 275836 334704 275888 334756
rect 278780 334704 278832 334756
rect 279240 334704 279292 334756
rect 333060 334636 333112 334688
rect 333244 334636 333296 334688
rect 244556 334432 244608 334484
rect 256700 334092 256752 334144
rect 257252 334092 257304 334144
rect 336832 333888 336884 333940
rect 337292 333888 337344 333940
rect 336832 333752 336884 333804
rect 337384 333752 337436 333804
rect 262772 333727 262824 333736
rect 262772 333693 262781 333727
rect 262781 333693 262815 333727
rect 262815 333693 262824 333727
rect 262772 333684 262824 333693
rect 288624 333548 288676 333600
rect 289176 333548 289228 333600
rect 274916 333480 274968 333532
rect 275192 333480 275244 333532
rect 288900 333480 288952 333532
rect 289544 333480 289596 333532
rect 261116 333276 261168 333328
rect 261392 333276 261444 333328
rect 293960 333276 294012 333328
rect 295064 333276 295116 333328
rect 306748 333276 306800 333328
rect 307484 333276 307536 333328
rect 261392 333140 261444 333192
rect 261852 333140 261904 333192
rect 294236 333140 294288 333192
rect 294420 333140 294472 333192
rect 308128 332936 308180 332988
rect 308864 332936 308916 332988
rect 298100 332732 298152 332784
rect 298744 332732 298796 332784
rect 236736 332664 236788 332716
rect 237196 332664 237248 332716
rect 283012 332664 283064 332716
rect 283472 332664 283524 332716
rect 263876 332324 263928 332376
rect 264704 332324 264756 332376
rect 326068 332256 326120 332308
rect 326804 332256 326856 332308
rect 246212 332052 246264 332104
rect 246672 332052 246724 332104
rect 287336 332052 287388 332104
rect 287888 332052 287940 332104
rect 241888 331984 241940 332036
rect 242164 331984 242216 332036
rect 231032 331848 231084 331900
rect 231308 331848 231360 331900
rect 272248 331848 272300 331900
rect 273076 331848 273128 331900
rect 311256 331848 311308 331900
rect 311440 331848 311492 331900
rect 329012 331848 329064 331900
rect 329564 331848 329616 331900
rect 333244 331848 333296 331900
rect 333704 331848 333756 331900
rect 323400 331712 323452 331764
rect 323860 331712 323912 331764
rect 298192 331372 298244 331424
rect 298836 331372 298888 331424
rect 301228 331304 301280 331356
rect 240784 331236 240836 331288
rect 245844 331236 245896 331288
rect 260196 331236 260248 331288
rect 260012 331168 260064 331220
rect 246028 331100 246080 331152
rect 298744 331100 298796 331152
rect 299204 331100 299256 331152
rect 304724 331236 304776 331288
rect 309876 331236 309928 331288
rect 304264 331168 304316 331220
rect 309692 331168 309744 331220
rect 290096 331032 290148 331084
rect 290372 331032 290424 331084
rect 301228 331032 301280 331084
rect 240692 330964 240744 331016
rect 295616 330828 295668 330880
rect 296536 330828 296588 330880
rect 258264 330692 258316 330744
rect 259368 330692 259420 330744
rect 341524 330624 341576 330676
rect 342076 330624 342128 330676
rect 302332 330556 302384 330608
rect 303160 330556 303212 330608
rect 320364 330556 320416 330608
rect 321376 330556 321428 330608
rect 323216 330556 323268 330608
rect 324228 330556 324280 330608
rect 288624 330488 288676 330540
rect 289360 330488 289412 330540
rect 321836 330488 321888 330540
rect 322664 330488 322716 330540
rect 323124 330488 323176 330540
rect 324044 330488 324096 330540
rect 321652 330420 321704 330472
rect 322756 330420 322808 330472
rect 322940 330420 322992 330472
rect 323952 330420 324004 330472
rect 321560 330352 321612 330404
rect 322480 330352 322532 330404
rect 317512 330284 317564 330336
rect 318616 330284 318668 330336
rect 305000 329944 305052 329996
rect 305460 329944 305512 329996
rect 245936 329128 245988 329180
rect 246120 329128 246172 329180
rect 295432 328720 295484 328772
rect 296352 328720 296404 328772
rect 242532 328516 242584 328568
rect 286140 328516 286192 328568
rect 299848 328516 299900 328568
rect 300124 328516 300176 328568
rect 301044 328516 301096 328568
rect 301596 328516 301648 328568
rect 306656 328516 306708 328568
rect 307576 328516 307628 328568
rect 232136 328491 232188 328500
rect 232136 328457 232145 328491
rect 232145 328457 232179 328491
rect 232179 328457 232188 328491
rect 232136 328448 232188 328457
rect 242256 328448 242308 328500
rect 243636 328448 243688 328500
rect 243820 328448 243872 328500
rect 244464 328491 244516 328500
rect 244464 328457 244473 328491
rect 244473 328457 244507 328491
rect 244507 328457 244516 328491
rect 244464 328448 244516 328457
rect 253112 328448 253164 328500
rect 253664 328448 253716 328500
rect 265440 328448 265492 328500
rect 265532 328448 265584 328500
rect 277584 328448 277636 328500
rect 278504 328448 278556 328500
rect 284668 328448 284720 328500
rect 285496 328448 285548 328500
rect 285864 328448 285916 328500
rect 285956 328448 286008 328500
rect 286600 328448 286652 328500
rect 326252 328448 326304 328500
rect 100668 328423 100720 328432
rect 100668 328389 100677 328423
rect 100677 328389 100711 328423
rect 100711 328389 100720 328423
rect 100668 328380 100720 328389
rect 231124 328423 231176 328432
rect 231124 328389 231133 328423
rect 231133 328389 231167 328423
rect 231167 328389 231176 328423
rect 231124 328380 231176 328389
rect 254676 328423 254728 328432
rect 254676 328389 254685 328423
rect 254685 328389 254719 328423
rect 254719 328389 254728 328423
rect 254676 328380 254728 328389
rect 258632 328380 258684 328432
rect 258816 328380 258868 328432
rect 263692 328380 263744 328432
rect 280620 328423 280672 328432
rect 280620 328389 280629 328423
rect 280629 328389 280663 328423
rect 280663 328389 280672 328423
rect 280620 328380 280672 328389
rect 281908 328423 281960 328432
rect 281908 328389 281917 328423
rect 281917 328389 281951 328423
rect 281951 328389 281960 328423
rect 281908 328380 281960 328389
rect 290280 328380 290332 328432
rect 290648 328380 290700 328432
rect 291752 328380 291804 328432
rect 291936 328380 291988 328432
rect 319444 328423 319496 328432
rect 319444 328389 319453 328423
rect 319453 328389 319487 328423
rect 319487 328389 319496 328423
rect 319444 328380 319496 328389
rect 326344 328380 326396 328432
rect 341524 328380 341576 328432
rect 341708 328380 341760 328432
rect 344284 328423 344336 328432
rect 344284 328389 344293 328423
rect 344293 328389 344327 328423
rect 344327 328389 344336 328423
rect 344284 328380 344336 328389
rect 263784 328312 263836 328364
rect 270500 328312 270552 328364
rect 271512 328312 271564 328364
rect 284484 328244 284536 328296
rect 285312 328244 285364 328296
rect 265256 328176 265308 328228
rect 266084 328176 266136 328228
rect 269580 327904 269632 327956
rect 270040 327904 270092 327956
rect 273628 327428 273680 327480
rect 274180 327428 274232 327480
rect 267832 327292 267884 327344
rect 268844 327292 268896 327344
rect 273444 327224 273496 327276
rect 273904 327224 273956 327276
rect 336188 327156 336240 327208
rect 107476 327131 107528 327140
rect 107476 327097 107485 327131
rect 107485 327097 107519 327131
rect 107519 327097 107528 327131
rect 107476 327088 107528 327097
rect 266820 327088 266872 327140
rect 267464 327088 267516 327140
rect 272340 327088 272392 327140
rect 272524 327088 272576 327140
rect 279516 327131 279568 327140
rect 279516 327097 279525 327131
rect 279525 327097 279559 327131
rect 279559 327097 279568 327131
rect 279516 327088 279568 327097
rect 334532 327088 334584 327140
rect 335176 327088 335228 327140
rect 335820 327088 335872 327140
rect 257068 327063 257120 327072
rect 257068 327029 257077 327063
rect 257077 327029 257111 327063
rect 257111 327029 257120 327063
rect 257068 327020 257120 327029
rect 295616 327063 295668 327072
rect 295616 327029 295625 327063
rect 295625 327029 295659 327063
rect 295659 327029 295668 327063
rect 295616 327020 295668 327029
rect 341708 327020 341760 327072
rect 287428 326952 287480 327004
rect 288072 326952 288124 327004
rect 270592 326680 270644 326732
rect 271604 326680 271656 326732
rect 270776 326612 270828 326664
rect 271420 326612 271472 326664
rect 297180 326544 297232 326596
rect 297916 326544 297968 326596
rect 262404 326476 262456 326528
rect 263324 326476 263376 326528
rect 282920 326476 282972 326528
rect 284116 326476 284168 326528
rect 289912 326476 289964 326528
rect 291108 326476 291160 326528
rect 291292 326476 291344 326528
rect 292488 326476 292540 326528
rect 292764 326476 292816 326528
rect 293776 326476 293828 326528
rect 297364 326476 297416 326528
rect 298008 326476 298060 326528
rect 307852 326476 307904 326528
rect 308956 326476 309008 326528
rect 311900 326476 311952 326528
rect 313096 326476 313148 326528
rect 313280 326476 313332 326528
rect 314568 326476 314620 326528
rect 315212 326476 315264 326528
rect 315856 326476 315908 326528
rect 318800 326476 318852 326528
rect 320088 326476 320140 326528
rect 259460 326408 259512 326460
rect 260564 326408 260616 326460
rect 260840 326408 260892 326460
rect 261852 326408 261904 326460
rect 262588 326408 262640 326460
rect 263416 326408 263468 326460
rect 264980 326408 265032 326460
rect 265900 326408 265952 326460
rect 266360 326408 266412 326460
rect 267372 326408 267424 326460
rect 267740 326408 267792 326460
rect 268936 326408 268988 326460
rect 269212 326408 269264 326460
rect 270316 326408 270368 326460
rect 273444 326408 273496 326460
rect 274272 326408 274324 326460
rect 275100 326408 275152 326460
rect 275928 326408 275980 326460
rect 276296 326408 276348 326460
rect 277032 326408 277084 326460
rect 277768 326408 277820 326460
rect 278688 326408 278740 326460
rect 278780 326408 278832 326460
rect 279884 326408 279936 326460
rect 280252 326408 280304 326460
rect 281448 326408 281500 326460
rect 281632 326408 281684 326460
rect 282552 326408 282604 326460
rect 283288 326408 283340 326460
rect 284024 326408 284076 326460
rect 284392 326408 284444 326460
rect 285588 326408 285640 326460
rect 285680 326408 285732 326460
rect 286968 326408 287020 326460
rect 287704 326408 287756 326460
rect 288348 326408 288400 326460
rect 288808 326408 288860 326460
rect 289544 326408 289596 326460
rect 290096 326408 290148 326460
rect 290924 326408 290976 326460
rect 291476 326408 291528 326460
rect 292212 326408 292264 326460
rect 292948 326408 293000 326460
rect 293592 326408 293644 326460
rect 294052 326408 294104 326460
rect 295248 326408 295300 326460
rect 295892 326408 295944 326460
rect 296536 326408 296588 326460
rect 298192 326408 298244 326460
rect 299388 326408 299440 326460
rect 301228 326408 301280 326460
rect 302148 326408 302200 326460
rect 302240 326408 302292 326460
rect 303436 326408 303488 326460
rect 304080 326408 304132 326460
rect 304816 326408 304868 326460
rect 305184 326408 305236 326460
rect 306196 326408 306248 326460
rect 306472 326408 306524 326460
rect 307668 326408 307720 326460
rect 308036 326408 308088 326460
rect 308864 326408 308916 326460
rect 309140 326408 309192 326460
rect 310244 326408 310296 326460
rect 311256 326408 311308 326460
rect 311716 326408 311768 326460
rect 312084 326408 312136 326460
rect 312820 326408 312872 326460
rect 313556 326408 313608 326460
rect 314384 326408 314436 326460
rect 317972 326408 318024 326460
rect 318432 326408 318484 326460
rect 319076 326408 319128 326460
rect 319812 326408 319864 326460
rect 258724 326340 258776 326392
rect 259276 326340 259328 326392
rect 259736 326340 259788 326392
rect 260748 326340 260800 326392
rect 261208 326340 261260 326392
rect 262036 326340 262088 326392
rect 262680 326340 262732 326392
rect 263232 326340 263284 326392
rect 263600 326340 263652 326392
rect 264796 326340 264848 326392
rect 265072 326340 265124 326392
rect 265992 326340 266044 326392
rect 266636 326340 266688 326392
rect 267556 326340 267608 326392
rect 268016 326340 268068 326392
rect 268752 326340 268804 326392
rect 270684 326340 270736 326392
rect 271788 326340 271840 326392
rect 271880 326340 271932 326392
rect 272984 326340 273036 326392
rect 273720 326340 273772 326392
rect 274364 326340 274416 326392
rect 274732 326340 274784 326392
rect 275652 326340 275704 326392
rect 276664 326340 276716 326392
rect 277216 326340 277268 326392
rect 277676 326340 277728 326392
rect 278596 326340 278648 326392
rect 278872 326340 278924 326392
rect 279792 326340 279844 326392
rect 280344 326340 280396 326392
rect 281172 326340 281224 326392
rect 281724 326340 281776 326392
rect 282460 326340 282512 326392
rect 283196 326340 283248 326392
rect 283932 326340 283984 326392
rect 284300 326340 284352 326392
rect 285496 326340 285548 326392
rect 285772 326340 285824 326392
rect 286876 326340 286928 326392
rect 287612 326340 287664 326392
rect 288164 326340 288216 326392
rect 288900 326340 288952 326392
rect 289452 326340 289504 326392
rect 290188 326340 290240 326392
rect 291016 326340 291068 326392
rect 291568 326340 291620 326392
rect 292120 326340 292172 326392
rect 293040 326340 293092 326392
rect 293500 326340 293552 326392
rect 294236 326340 294288 326392
rect 295064 326340 295116 326392
rect 295340 326340 295392 326392
rect 296628 326340 296680 326392
rect 296720 326340 296772 326392
rect 297732 326340 297784 326392
rect 298376 326340 298428 326392
rect 299296 326340 299348 326392
rect 302700 326340 302752 326392
rect 303528 326340 303580 326392
rect 303804 326340 303856 326392
rect 304632 326340 304684 326392
rect 305092 326340 305144 326392
rect 306104 326340 306156 326392
rect 306564 326340 306616 326392
rect 307484 326340 307536 326392
rect 308128 326340 308180 326392
rect 308680 326340 308732 326392
rect 310612 326340 310664 326392
rect 311808 326340 311860 326392
rect 312360 326340 312412 326392
rect 312912 326340 312964 326392
rect 313648 326340 313700 326392
rect 314292 326340 314344 326392
rect 314752 326340 314804 326392
rect 315948 326340 316000 326392
rect 316224 326340 316276 326392
rect 317236 326340 317288 326392
rect 318064 326340 318116 326392
rect 318524 326340 318576 326392
rect 319168 326340 319220 326392
rect 319720 326340 319772 326392
rect 320456 326340 320508 326392
rect 321284 326340 321336 326392
rect 260932 326272 260984 326324
rect 262128 326272 262180 326324
rect 262220 326272 262272 326324
rect 263140 326272 263192 326324
rect 265164 326272 265216 326324
rect 266176 326272 266228 326324
rect 266544 326272 266596 326324
rect 267648 326272 267700 326324
rect 273260 326272 273312 326324
rect 274548 326272 274600 326324
rect 276112 326272 276164 326324
rect 276940 326272 276992 326324
rect 277400 326272 277452 326324
rect 278320 326272 278372 326324
rect 279056 326272 279108 326324
rect 280068 326272 280120 326324
rect 281540 326272 281592 326324
rect 282736 326272 282788 326324
rect 283012 326272 283064 326324
rect 284208 326272 284260 326324
rect 287336 326272 287388 326324
rect 288256 326272 288308 326324
rect 288440 326272 288492 326324
rect 289728 326272 289780 326324
rect 289820 326272 289872 326324
rect 290832 326272 290884 326324
rect 291660 326272 291712 326324
rect 292396 326272 292448 326324
rect 292856 326272 292908 326324
rect 293684 326272 293736 326324
rect 303620 326272 303672 326324
rect 304908 326272 304960 326324
rect 305000 326272 305052 326324
rect 306288 326272 306340 326324
rect 307944 326272 307996 326324
rect 308772 326272 308824 326324
rect 309232 326272 309284 326324
rect 310428 326272 310480 326324
rect 312176 326272 312228 326324
rect 313004 326272 313056 326324
rect 313372 326272 313424 326324
rect 314476 326272 314528 326324
rect 317696 326272 317748 326324
rect 318708 326272 318760 326324
rect 318984 326272 319036 326324
rect 319996 326272 320048 326324
rect 256976 326204 257028 326256
rect 257712 326204 257764 326256
rect 262496 326204 262548 326256
rect 263508 326204 263560 326256
rect 292580 326204 292632 326256
rect 293868 326204 293920 326256
rect 299664 326204 299716 326256
rect 300492 326204 300544 326256
rect 300860 326204 300912 326256
rect 301872 326204 301924 326256
rect 307760 326204 307812 326256
rect 309048 326204 309100 326256
rect 310704 326204 310756 326256
rect 311440 326204 311492 326256
rect 314844 326204 314896 326256
rect 315580 326204 315632 326256
rect 256792 326136 256844 326188
rect 257804 326136 257856 326188
rect 299480 326136 299532 326188
rect 300400 326136 300452 326188
rect 299572 326068 299624 326120
rect 300584 326068 300636 326120
rect 262864 325660 262916 325712
rect 318156 325660 318208 325712
rect 318248 325660 318300 325712
rect 319444 325703 319496 325712
rect 319444 325669 319453 325703
rect 319453 325669 319487 325703
rect 319487 325669 319496 325703
rect 319444 325660 319496 325669
rect 320272 325703 320324 325712
rect 320272 325669 320281 325703
rect 320281 325669 320315 325703
rect 320315 325669 320324 325703
rect 320272 325660 320324 325669
rect 330760 325660 330812 325712
rect 330944 325660 330996 325712
rect 335820 325635 335872 325644
rect 335820 325601 335829 325635
rect 335829 325601 335863 325635
rect 335863 325601 335872 325635
rect 335820 325592 335872 325601
rect 296904 325524 296956 325576
rect 297548 325524 297600 325576
rect 272248 324912 272300 324964
rect 272800 324912 272852 324964
rect 268108 324708 268160 324760
rect 268660 324708 268712 324760
rect 261116 324436 261168 324488
rect 261576 324436 261628 324488
rect 2780 324164 2832 324216
rect 4712 324164 4764 324216
rect 275008 323552 275060 323604
rect 275560 323552 275612 323604
rect 298468 323552 298520 323604
rect 299112 323552 299164 323604
rect 305460 323552 305512 323604
rect 305920 323552 305972 323604
rect 309508 323552 309560 323604
rect 310336 323552 310388 323604
rect 298100 323416 298152 323468
rect 299020 323416 299072 323468
rect 262864 322192 262916 322244
rect 263048 322192 263100 322244
rect 296076 322192 296128 322244
rect 244464 321580 244516 321632
rect 259736 321512 259788 321564
rect 260380 321512 260432 321564
rect 309416 321512 309468 321564
rect 310060 321512 310112 321564
rect 310888 321512 310940 321564
rect 311348 321512 311400 321564
rect 244464 321444 244516 321496
rect 266912 321444 266964 321496
rect 267188 321444 267240 321496
rect 277584 321444 277636 321496
rect 278228 321444 278280 321496
rect 302608 321444 302660 321496
rect 303068 321444 303120 321496
rect 303896 321444 303948 321496
rect 304448 321444 304500 321496
rect 100668 318835 100720 318844
rect 100668 318801 100677 318835
rect 100677 318801 100711 318835
rect 100711 318801 100720 318835
rect 100668 318792 100720 318801
rect 231216 318792 231268 318844
rect 232320 318792 232372 318844
rect 232412 318792 232464 318844
rect 232596 318792 232648 318844
rect 232688 318792 232740 318844
rect 254860 318792 254912 318844
rect 265624 318792 265676 318844
rect 272524 318792 272576 318844
rect 272892 318792 272944 318844
rect 273812 318792 273864 318844
rect 274088 318792 274140 318844
rect 280988 318792 281040 318844
rect 282368 318792 282420 318844
rect 344376 318792 344428 318844
rect 315028 318724 315080 318776
rect 315488 318724 315540 318776
rect 265808 318656 265860 318708
rect 282644 318699 282696 318708
rect 282644 318665 282653 318699
rect 282653 318665 282687 318699
rect 282687 318665 282696 318699
rect 282644 318656 282696 318665
rect 258724 317500 258776 317552
rect 258908 317500 258960 317552
rect 257160 317432 257212 317484
rect 293316 317432 293368 317484
rect 293408 317432 293460 317484
rect 293960 317432 294012 317484
rect 294788 317432 294840 317484
rect 341616 317475 341668 317484
rect 341616 317441 341625 317475
rect 341625 317441 341659 317475
rect 341659 317441 341668 317475
rect 341616 317432 341668 317441
rect 107476 317407 107528 317416
rect 107476 317373 107485 317407
rect 107485 317373 107519 317407
rect 107519 317373 107528 317407
rect 107476 317364 107528 317373
rect 232320 317364 232372 317416
rect 232412 317364 232464 317416
rect 244372 317407 244424 317416
rect 244372 317373 244381 317407
rect 244381 317373 244415 317407
rect 244415 317373 244424 317407
rect 244372 317364 244424 317373
rect 260380 317407 260432 317416
rect 260380 317373 260389 317407
rect 260389 317373 260423 317407
rect 260423 317373 260432 317407
rect 260380 317364 260432 317373
rect 261668 317364 261720 317416
rect 265808 317407 265860 317416
rect 265808 317373 265817 317407
rect 265817 317373 265851 317407
rect 265851 317373 265860 317407
rect 265808 317364 265860 317373
rect 331772 317364 331824 317416
rect 331864 317364 331916 317416
rect 333060 317364 333112 317416
rect 333152 317364 333204 317416
rect 333244 317364 333296 317416
rect 333336 317364 333388 317416
rect 340144 317364 340196 317416
rect 271972 316684 272024 316736
rect 272708 316684 272760 316736
rect 284576 316548 284628 316600
rect 316132 316548 316184 316600
rect 316868 316548 316920 316600
rect 285036 316480 285088 316532
rect 319444 316072 319496 316124
rect 319628 316072 319680 316124
rect 301044 316004 301096 316056
rect 301780 316004 301832 316056
rect 330576 316004 330628 316056
rect 330760 316004 330812 316056
rect 336004 316004 336056 316056
rect 258908 315936 258960 315988
rect 319444 315979 319496 315988
rect 319444 315945 319453 315979
rect 319453 315945 319487 315979
rect 319487 315945 319496 315979
rect 319444 315936 319496 315945
rect 320272 315979 320324 315988
rect 320272 315945 320281 315979
rect 320281 315945 320315 315979
rect 320315 315945 320324 315979
rect 320272 315936 320324 315945
rect 317880 315188 317932 315240
rect 318248 315188 318300 315240
rect 285864 313896 285916 313948
rect 286508 313896 286560 313948
rect 263784 313488 263836 313540
rect 264520 313488 264572 313540
rect 322296 312672 322348 312724
rect 322572 312672 322624 312724
rect 231216 311924 231268 311976
rect 289268 311924 289320 311976
rect 344192 311856 344244 311908
rect 344376 311856 344428 311908
rect 289176 311788 289228 311840
rect 231216 311720 231268 311772
rect 244372 311491 244424 311500
rect 244372 311457 244381 311491
rect 244381 311457 244415 311491
rect 244415 311457 244424 311491
rect 244372 311448 244424 311457
rect 322296 311108 322348 311160
rect 322572 311108 322624 311160
rect 310060 309884 310112 309936
rect 311348 309884 311400 309936
rect 310060 309748 310112 309800
rect 311348 309748 311400 309800
rect 280896 309136 280948 309188
rect 280988 309136 281040 309188
rect 282644 309179 282696 309188
rect 282644 309145 282653 309179
rect 282653 309145 282687 309179
rect 282687 309145 282696 309179
rect 282644 309136 282696 309145
rect 293316 309136 293368 309188
rect 100668 309111 100720 309120
rect 100668 309077 100677 309111
rect 100677 309077 100711 309111
rect 100711 309077 100720 309111
rect 100668 309068 100720 309077
rect 238024 309111 238076 309120
rect 238024 309077 238033 309111
rect 238033 309077 238067 309111
rect 238067 309077 238076 309111
rect 238024 309068 238076 309077
rect 246396 309068 246448 309120
rect 253112 309068 253164 309120
rect 253204 309068 253256 309120
rect 254676 309068 254728 309120
rect 254860 309068 254912 309120
rect 257068 309068 257120 309120
rect 257160 309068 257212 309120
rect 326252 309068 326304 309120
rect 326344 309068 326396 309120
rect 246488 309000 246540 309052
rect 265808 307887 265860 307896
rect 265808 307853 265817 307887
rect 265817 307853 265851 307887
rect 265851 307853 265860 307887
rect 265808 307844 265860 307853
rect 107476 307819 107528 307828
rect 107476 307785 107485 307819
rect 107485 307785 107519 307819
rect 107519 307785 107528 307819
rect 107476 307776 107528 307785
rect 260380 307819 260432 307828
rect 260380 307785 260389 307819
rect 260389 307785 260423 307819
rect 260423 307785 260432 307819
rect 260380 307776 260432 307785
rect 329012 307776 329064 307828
rect 329104 307776 329156 307828
rect 339960 307819 340012 307828
rect 339960 307785 339969 307819
rect 339969 307785 340003 307819
rect 340003 307785 340012 307819
rect 339960 307776 340012 307785
rect 264520 307751 264572 307760
rect 264520 307717 264529 307751
rect 264529 307717 264563 307751
rect 264563 307717 264572 307751
rect 264520 307708 264572 307717
rect 265808 307751 265860 307760
rect 265808 307717 265817 307751
rect 265817 307717 265851 307751
rect 265851 307717 265860 307751
rect 265808 307708 265860 307717
rect 316868 307751 316920 307760
rect 316868 307717 316877 307751
rect 316877 307717 316911 307751
rect 316911 307717 316920 307751
rect 316868 307708 316920 307717
rect 318064 307028 318116 307080
rect 318340 307028 318392 307080
rect 293408 306391 293460 306400
rect 293408 306357 293417 306391
rect 293417 306357 293451 306391
rect 293451 306357 293460 306391
rect 293408 306348 293460 306357
rect 319628 306348 319680 306400
rect 321100 306348 321152 306400
rect 335820 306348 335872 306400
rect 336004 306348 336056 306400
rect 267188 304308 267240 304360
rect 268660 304308 268712 304360
rect 267188 304172 267240 304224
rect 268660 304172 268712 304224
rect 257068 302923 257120 302932
rect 257068 302889 257077 302923
rect 257077 302889 257111 302923
rect 257111 302889 257120 302923
rect 257068 302880 257120 302889
rect 341616 302200 341668 302252
rect 341708 302064 341760 302116
rect 100668 299523 100720 299532
rect 100668 299489 100677 299523
rect 100677 299489 100711 299523
rect 100711 299489 100720 299523
rect 100668 299480 100720 299489
rect 238024 299523 238076 299532
rect 238024 299489 238033 299523
rect 238033 299489 238067 299523
rect 238067 299489 238076 299523
rect 238024 299480 238076 299489
rect 244924 299480 244976 299532
rect 245016 299480 245068 299532
rect 254676 299480 254728 299532
rect 261576 299523 261628 299532
rect 261576 299489 261585 299523
rect 261585 299489 261619 299523
rect 261619 299489 261628 299523
rect 261576 299480 261628 299489
rect 322204 299480 322256 299532
rect 322296 299480 322348 299532
rect 231216 299455 231268 299464
rect 231216 299421 231225 299455
rect 231225 299421 231259 299455
rect 231259 299421 231268 299455
rect 231216 299412 231268 299421
rect 231952 299412 232004 299464
rect 232044 299412 232096 299464
rect 232320 299412 232372 299464
rect 232412 299412 232464 299464
rect 240692 299455 240744 299464
rect 240692 299421 240701 299455
rect 240701 299421 240735 299455
rect 240735 299421 240744 299455
rect 240692 299412 240744 299421
rect 246396 299412 246448 299464
rect 246488 299412 246540 299464
rect 260288 299455 260340 299464
rect 260288 299421 260297 299455
rect 260297 299421 260331 299455
rect 260331 299421 260340 299455
rect 260288 299412 260340 299421
rect 331772 299412 331824 299464
rect 331864 299412 331916 299464
rect 333244 299412 333296 299464
rect 333336 299412 333388 299464
rect 334532 299412 334584 299464
rect 334624 299412 334676 299464
rect 339960 299412 340012 299464
rect 340144 299412 340196 299464
rect 341708 299412 341760 299464
rect 345388 299412 345440 299464
rect 254860 299344 254912 299396
rect 341708 299276 341760 299328
rect 345388 299276 345440 299328
rect 258816 298163 258868 298172
rect 258816 298129 258825 298163
rect 258825 298129 258859 298163
rect 258859 298129 258868 298163
rect 258816 298120 258868 298129
rect 264520 298163 264572 298172
rect 264520 298129 264529 298163
rect 264529 298129 264563 298163
rect 264563 298129 264572 298163
rect 264520 298120 264572 298129
rect 265808 298163 265860 298172
rect 265808 298129 265817 298163
rect 265817 298129 265851 298163
rect 265851 298129 265860 298163
rect 265808 298120 265860 298129
rect 293316 298120 293368 298172
rect 293408 298120 293460 298172
rect 316960 298120 317012 298172
rect 107476 298095 107528 298104
rect 107476 298061 107485 298095
rect 107485 298061 107519 298095
rect 107519 298061 107528 298095
rect 107476 298052 107528 298061
rect 231952 298052 232004 298104
rect 232044 298052 232096 298104
rect 232412 298095 232464 298104
rect 232412 298061 232421 298095
rect 232421 298061 232455 298095
rect 232455 298061 232464 298095
rect 232412 298052 232464 298061
rect 245016 298095 245068 298104
rect 245016 298061 245025 298095
rect 245025 298061 245059 298095
rect 245059 298061 245068 298095
rect 245016 298052 245068 298061
rect 319628 298095 319680 298104
rect 319628 298061 319637 298095
rect 319637 298061 319671 298095
rect 319671 298061 319680 298095
rect 319628 298052 319680 298061
rect 321100 298095 321152 298104
rect 321100 298061 321109 298095
rect 321109 298061 321143 298095
rect 321143 298061 321152 298095
rect 321100 298052 321152 298061
rect 333244 298052 333296 298104
rect 333336 298052 333388 298104
rect 339960 298095 340012 298104
rect 339960 298061 339969 298095
rect 339969 298061 340003 298095
rect 340003 298061 340012 298095
rect 339960 298052 340012 298061
rect 335912 296692 335964 296744
rect 336004 296692 336056 296744
rect 257160 294448 257212 294500
rect 232688 292612 232740 292664
rect 232688 292476 232740 292528
rect 333152 290003 333204 290012
rect 333152 289969 333161 290003
rect 333161 289969 333195 290003
rect 333195 289969 333204 290003
rect 333152 289960 333204 289969
rect 231216 289867 231268 289876
rect 231216 289833 231225 289867
rect 231225 289833 231259 289867
rect 231259 289833 231268 289867
rect 231216 289824 231268 289833
rect 240692 289867 240744 289876
rect 240692 289833 240701 289867
rect 240701 289833 240735 289867
rect 240735 289833 240744 289867
rect 240692 289824 240744 289833
rect 244372 289824 244424 289876
rect 244464 289824 244516 289876
rect 253020 289824 253072 289876
rect 253204 289824 253256 289876
rect 260380 289824 260432 289876
rect 322204 289824 322256 289876
rect 100668 289799 100720 289808
rect 100668 289765 100677 289799
rect 100677 289765 100711 289799
rect 100711 289765 100720 289799
rect 100668 289756 100720 289765
rect 238024 289799 238076 289808
rect 238024 289765 238033 289799
rect 238033 289765 238067 289799
rect 238067 289765 238076 289799
rect 238024 289756 238076 289765
rect 261484 289756 261536 289808
rect 261576 289756 261628 289808
rect 331864 289824 331916 289876
rect 334624 289824 334676 289876
rect 331772 289756 331824 289808
rect 334532 289756 334584 289808
rect 322204 289688 322256 289740
rect 321100 288507 321152 288516
rect 321100 288473 321109 288507
rect 321109 288473 321143 288507
rect 321143 288473 321152 288507
rect 321100 288464 321152 288473
rect 329012 288464 329064 288516
rect 329196 288464 329248 288516
rect 330576 288464 330628 288516
rect 335820 288464 335872 288516
rect 336004 288464 336056 288516
rect 107476 288439 107528 288448
rect 107476 288405 107485 288439
rect 107485 288405 107519 288439
rect 107519 288405 107528 288439
rect 107476 288396 107528 288405
rect 232412 288439 232464 288448
rect 232412 288405 232421 288439
rect 232421 288405 232455 288439
rect 232455 288405 232464 288439
rect 232412 288396 232464 288405
rect 254860 288396 254912 288448
rect 254952 288396 255004 288448
rect 293224 288396 293276 288448
rect 293316 288396 293368 288448
rect 330484 288396 330536 288448
rect 333152 288439 333204 288448
rect 333152 288405 333161 288439
rect 333161 288405 333195 288439
rect 333195 288405 333204 288439
rect 333152 288396 333204 288405
rect 246396 288371 246448 288380
rect 246396 288337 246405 288371
rect 246405 288337 246439 288371
rect 246439 288337 246448 288371
rect 246396 288328 246448 288337
rect 265808 288371 265860 288380
rect 265808 288337 265817 288371
rect 265817 288337 265851 288371
rect 265851 288337 265860 288371
rect 265808 288328 265860 288337
rect 319628 287079 319680 287088
rect 319628 287045 319637 287079
rect 319637 287045 319671 287079
rect 319671 287045 319680 287079
rect 319628 287036 319680 287045
rect 326252 287036 326304 287088
rect 326436 287036 326488 287088
rect 258908 286968 258960 287020
rect 340052 282820 340104 282872
rect 100668 280211 100720 280220
rect 100668 280177 100677 280211
rect 100677 280177 100711 280211
rect 100711 280177 100720 280211
rect 100668 280168 100720 280177
rect 238024 280211 238076 280220
rect 238024 280177 238033 280211
rect 238033 280177 238067 280211
rect 238067 280177 238076 280211
rect 238024 280168 238076 280177
rect 254768 280168 254820 280220
rect 254860 280168 254912 280220
rect 2780 280100 2832 280152
rect 5448 280100 5500 280152
rect 231216 280143 231268 280152
rect 231216 280109 231225 280143
rect 231225 280109 231259 280143
rect 231259 280109 231268 280143
rect 231216 280100 231268 280109
rect 232044 280100 232096 280152
rect 232136 280100 232188 280152
rect 240692 280143 240744 280152
rect 240692 280109 240701 280143
rect 240701 280109 240735 280143
rect 240735 280109 240744 280143
rect 240692 280100 240744 280109
rect 246028 280143 246080 280152
rect 246028 280109 246037 280143
rect 246037 280109 246071 280143
rect 246071 280109 246080 280143
rect 246028 280100 246080 280109
rect 257160 280143 257212 280152
rect 257160 280109 257169 280143
rect 257169 280109 257203 280143
rect 257203 280109 257212 280143
rect 257160 280100 257212 280109
rect 330484 280100 330536 280152
rect 330576 280100 330628 280152
rect 331772 280100 331824 280152
rect 331864 280100 331916 280152
rect 333244 280100 333296 280152
rect 333336 280100 333388 280152
rect 334532 280100 334584 280152
rect 334624 280100 334676 280152
rect 340052 280100 340104 280152
rect 340144 280100 340196 280152
rect 265808 278851 265860 278860
rect 265808 278817 265817 278851
rect 265817 278817 265851 278851
rect 265851 278817 265860 278851
rect 265808 278808 265860 278817
rect 244464 278740 244516 278792
rect 244648 278740 244700 278792
rect 244924 278740 244976 278792
rect 246488 278740 246540 278792
rect 257160 278783 257212 278792
rect 257160 278749 257169 278783
rect 257169 278749 257203 278783
rect 257203 278749 257212 278783
rect 257160 278740 257212 278749
rect 293132 278740 293184 278792
rect 293316 278740 293368 278792
rect 329012 278740 329064 278792
rect 329196 278740 329248 278792
rect 335820 278740 335872 278792
rect 336004 278740 336056 278792
rect 264520 278715 264572 278724
rect 264520 278681 264529 278715
rect 264529 278681 264563 278715
rect 264563 278681 264572 278715
rect 264520 278672 264572 278681
rect 265808 278715 265860 278724
rect 265808 278681 265817 278715
rect 265817 278681 265851 278715
rect 265851 278681 265860 278715
rect 265808 278672 265860 278681
rect 258724 277423 258776 277432
rect 258724 277389 258733 277423
rect 258733 277389 258767 277423
rect 258767 277389 258776 277423
rect 258724 277380 258776 277389
rect 232688 273300 232740 273352
rect 341616 273300 341668 273352
rect 260288 273275 260340 273284
rect 260288 273241 260297 273275
rect 260297 273241 260331 273275
rect 260331 273241 260340 273275
rect 260288 273232 260340 273241
rect 333152 273232 333204 273284
rect 232688 273164 232740 273216
rect 333060 273164 333112 273216
rect 341616 273164 341668 273216
rect 246488 272552 246540 272604
rect 246764 272552 246816 272604
rect 328920 270580 328972 270632
rect 231216 270555 231268 270564
rect 231216 270521 231225 270555
rect 231225 270521 231259 270555
rect 231259 270521 231268 270555
rect 231216 270512 231268 270521
rect 240692 270555 240744 270564
rect 240692 270521 240701 270555
rect 240701 270521 240735 270555
rect 240735 270521 240744 270555
rect 240692 270512 240744 270521
rect 246028 270555 246080 270564
rect 246028 270521 246037 270555
rect 246037 270521 246071 270555
rect 246071 270521 246080 270555
rect 246028 270512 246080 270521
rect 345296 270512 345348 270564
rect 345388 270512 345440 270564
rect 100668 270487 100720 270496
rect 100668 270453 100677 270487
rect 100677 270453 100711 270487
rect 100711 270453 100720 270487
rect 100668 270444 100720 270453
rect 238024 270487 238076 270496
rect 238024 270453 238033 270487
rect 238033 270453 238067 270487
rect 238067 270453 238076 270487
rect 238024 270444 238076 270453
rect 244924 270444 244976 270496
rect 245108 270444 245160 270496
rect 328920 270444 328972 270496
rect 107476 269084 107528 269136
rect 107660 269084 107712 269136
rect 231952 269084 232004 269136
rect 232136 269084 232188 269136
rect 261392 269084 261444 269136
rect 261668 269084 261720 269136
rect 264520 269127 264572 269136
rect 264520 269093 264529 269127
rect 264529 269093 264563 269127
rect 264563 269093 264572 269127
rect 264520 269084 264572 269093
rect 265808 269127 265860 269136
rect 265808 269093 265817 269127
rect 265817 269093 265851 269127
rect 265851 269093 265860 269127
rect 265808 269084 265860 269093
rect 320916 269084 320968 269136
rect 321100 269084 321152 269136
rect 319444 267724 319496 267776
rect 319628 267724 319680 267776
rect 326344 267724 326396 267776
rect 326528 267724 326580 267776
rect 331588 266296 331640 266348
rect 331864 266296 331916 266348
rect 2780 266092 2832 266144
rect 5356 266092 5408 266144
rect 260380 265276 260432 265328
rect 322296 263619 322348 263628
rect 322296 263585 322305 263619
rect 322305 263585 322339 263619
rect 322339 263585 322348 263619
rect 322296 263576 322348 263585
rect 333060 263576 333112 263628
rect 333152 263508 333204 263560
rect 231768 262896 231820 262948
rect 232044 262896 232096 262948
rect 100668 260899 100720 260908
rect 100668 260865 100677 260899
rect 100677 260865 100711 260899
rect 100711 260865 100720 260899
rect 100668 260856 100720 260865
rect 238024 260899 238076 260908
rect 238024 260865 238033 260899
rect 238033 260865 238067 260899
rect 238067 260865 238076 260899
rect 238024 260856 238076 260865
rect 328920 260856 328972 260908
rect 329012 260856 329064 260908
rect 333244 260856 333296 260908
rect 333336 260856 333388 260908
rect 334532 260856 334584 260908
rect 334624 260856 334676 260908
rect 335728 260856 335780 260908
rect 335820 260856 335872 260908
rect 231216 260831 231268 260840
rect 231216 260797 231225 260831
rect 231225 260797 231259 260831
rect 231259 260797 231268 260831
rect 231216 260788 231268 260797
rect 330484 260788 330536 260840
rect 330576 260788 330628 260840
rect 341616 260831 341668 260840
rect 341616 260797 341625 260831
rect 341625 260797 341659 260831
rect 341659 260797 341668 260831
rect 341616 260788 341668 260797
rect 345388 260788 345440 260840
rect 345388 260652 345440 260704
rect 257068 259428 257120 259480
rect 257160 259428 257212 259480
rect 264336 259428 264388 259480
rect 264520 259428 264572 259480
rect 265624 259428 265676 259480
rect 265808 259428 265860 259480
rect 293132 259428 293184 259480
rect 293316 259428 293368 259480
rect 320916 259428 320968 259480
rect 321100 259428 321152 259480
rect 322296 259471 322348 259480
rect 322296 259437 322305 259471
rect 322305 259437 322339 259471
rect 322339 259437 322348 259471
rect 322296 259428 322348 259437
rect 244924 259360 244976 259412
rect 245108 259360 245160 259412
rect 246304 258068 246356 258120
rect 246396 258068 246448 258120
rect 258632 258068 258684 258120
rect 258724 258068 258776 258120
rect 232044 258000 232096 258052
rect 232320 258000 232372 258052
rect 244372 258043 244424 258052
rect 244372 258009 244381 258043
rect 244381 258009 244415 258043
rect 244415 258009 244424 258043
rect 244372 258000 244424 258009
rect 319628 258043 319680 258052
rect 319628 258009 319637 258043
rect 319637 258009 319671 258043
rect 319671 258009 319680 258043
rect 319628 258000 319680 258009
rect 322112 258000 322164 258052
rect 322204 258000 322256 258052
rect 335820 258000 335872 258052
rect 299020 256683 299072 256692
rect 299020 256649 299029 256683
rect 299029 256649 299063 256683
rect 299063 256649 299072 256683
rect 299020 256640 299072 256649
rect 334532 256683 334584 256692
rect 334532 256649 334541 256683
rect 334541 256649 334575 256683
rect 334575 256649 334584 256683
rect 334532 256640 334584 256649
rect 326344 254056 326396 254108
rect 253112 253988 253164 254040
rect 333152 253920 333204 253972
rect 232136 253895 232188 253904
rect 232136 253861 232145 253895
rect 232145 253861 232179 253895
rect 232179 253861 232188 253895
rect 232136 253852 232188 253861
rect 253020 253852 253072 253904
rect 333060 253852 333112 253904
rect 232320 253172 232372 253224
rect 265624 253172 265676 253224
rect 265808 253172 265860 253224
rect 231216 251243 231268 251252
rect 231216 251209 231225 251243
rect 231225 251209 231259 251243
rect 231259 251209 231268 251243
rect 231216 251200 231268 251209
rect 256976 251243 257028 251252
rect 256976 251209 256985 251243
rect 256985 251209 257019 251243
rect 257019 251209 257028 251243
rect 256976 251200 257028 251209
rect 341708 251200 341760 251252
rect 100668 251175 100720 251184
rect 100668 251141 100677 251175
rect 100677 251141 100711 251175
rect 100711 251141 100720 251175
rect 100668 251132 100720 251141
rect 334532 251107 334584 251116
rect 334532 251073 334541 251107
rect 334541 251073 334575 251107
rect 334575 251073 334584 251107
rect 334532 251064 334584 251073
rect 335820 250928 335872 250980
rect 258632 249840 258684 249892
rect 107476 249772 107528 249824
rect 107660 249772 107712 249824
rect 256976 249815 257028 249824
rect 256976 249781 256985 249815
rect 256985 249781 257019 249815
rect 257019 249781 257028 249815
rect 256976 249772 257028 249781
rect 258724 249772 258776 249824
rect 320916 249772 320968 249824
rect 321100 249772 321152 249824
rect 326252 249815 326304 249824
rect 326252 249781 326261 249815
rect 326261 249781 326295 249815
rect 326295 249781 326304 249815
rect 326252 249772 326304 249781
rect 345388 249772 345440 249824
rect 345572 249772 345624 249824
rect 258816 249747 258868 249756
rect 258816 249713 258825 249747
rect 258825 249713 258859 249747
rect 258859 249713 258868 249747
rect 258816 249704 258868 249713
rect 246304 248387 246356 248396
rect 246304 248353 246313 248387
rect 246313 248353 246347 248387
rect 246347 248353 246356 248387
rect 246304 248344 246356 248353
rect 299020 247095 299072 247104
rect 299020 247061 299029 247095
rect 299029 247061 299063 247095
rect 299063 247061 299072 247095
rect 299020 247052 299072 247061
rect 300308 247027 300360 247036
rect 300308 246993 300317 247027
rect 300317 246993 300351 247027
rect 300351 246993 300360 247027
rect 300308 246984 300360 246993
rect 301780 247027 301832 247036
rect 301780 246993 301789 247027
rect 301789 246993 301823 247027
rect 301823 246993 301832 247027
rect 301780 246984 301832 246993
rect 330484 246984 330536 247036
rect 330576 246984 330628 247036
rect 331772 246984 331824 247036
rect 331956 246984 332008 247036
rect 333244 246984 333296 247036
rect 333428 246984 333480 247036
rect 333060 244264 333112 244316
rect 340052 244264 340104 244316
rect 344100 244264 344152 244316
rect 344284 244264 344336 244316
rect 333152 244196 333204 244248
rect 340144 244128 340196 244180
rect 244372 241587 244424 241596
rect 244372 241553 244381 241587
rect 244381 241553 244415 241587
rect 244415 241553 244424 241587
rect 244372 241544 244424 241553
rect 100668 241519 100720 241528
rect 100668 241485 100677 241519
rect 100677 241485 100711 241519
rect 100711 241485 100720 241519
rect 100668 241476 100720 241485
rect 253020 241476 253072 241528
rect 253112 241476 253164 241528
rect 335820 241476 335872 241528
rect 336004 241476 336056 241528
rect 260196 240252 260248 240304
rect 258816 240227 258868 240236
rect 258816 240193 258825 240227
rect 258825 240193 258859 240227
rect 258859 240193 258868 240227
rect 258816 240184 258868 240193
rect 232044 240116 232096 240168
rect 232136 240116 232188 240168
rect 260288 240116 260340 240168
rect 261484 240116 261536 240168
rect 261576 240116 261628 240168
rect 264336 240116 264388 240168
rect 264520 240116 264572 240168
rect 293132 240116 293184 240168
rect 293316 240116 293368 240168
rect 319628 240159 319680 240168
rect 319628 240125 319637 240159
rect 319637 240125 319671 240159
rect 319671 240125 319680 240159
rect 319628 240116 319680 240125
rect 320916 240116 320968 240168
rect 321100 240116 321152 240168
rect 232688 240091 232740 240100
rect 232688 240057 232697 240091
rect 232697 240057 232731 240091
rect 232731 240057 232740 240091
rect 232688 240048 232740 240057
rect 258632 240048 258684 240100
rect 258816 240048 258868 240100
rect 246396 238756 246448 238808
rect 261576 238731 261628 238740
rect 261576 238697 261585 238731
rect 261585 238697 261619 238731
rect 261619 238697 261628 238731
rect 261576 238688 261628 238697
rect 265624 238688 265676 238740
rect 265808 238688 265860 238740
rect 319444 238688 319496 238740
rect 319628 238688 319680 238740
rect 322112 238688 322164 238740
rect 322296 238688 322348 238740
rect 300308 237439 300360 237448
rect 300308 237405 300317 237439
rect 300317 237405 300351 237439
rect 300351 237405 300360 237439
rect 300308 237396 300360 237405
rect 301780 237439 301832 237448
rect 301780 237405 301789 237439
rect 301789 237405 301823 237439
rect 301823 237405 301832 237439
rect 301780 237396 301832 237405
rect 299020 237371 299072 237380
rect 299020 237337 299029 237371
rect 299029 237337 299063 237371
rect 299063 237337 299072 237371
rect 299020 237328 299072 237337
rect 329012 237328 329064 237380
rect 329196 237328 329248 237380
rect 330392 237328 330444 237380
rect 330484 237328 330536 237380
rect 2780 237260 2832 237312
rect 5264 237260 5316 237312
rect 301780 235943 301832 235952
rect 301780 235909 301789 235943
rect 301789 235909 301823 235943
rect 301823 235909 301832 235943
rect 301780 235900 301832 235909
rect 330392 235943 330444 235952
rect 330392 235909 330401 235943
rect 330401 235909 330435 235943
rect 330435 235909 330444 235943
rect 330392 235900 330444 235909
rect 232688 235331 232740 235340
rect 232688 235297 232697 235331
rect 232697 235297 232731 235331
rect 232731 235297 232740 235331
rect 232688 235288 232740 235297
rect 232044 234651 232096 234660
rect 232044 234617 232053 234651
rect 232053 234617 232087 234651
rect 232087 234617 232096 234651
rect 232044 234608 232096 234617
rect 245016 234608 245068 234660
rect 246396 234608 246448 234660
rect 244188 234540 244240 234592
rect 244372 234540 244424 234592
rect 244924 234540 244976 234592
rect 261576 234583 261628 234592
rect 261576 234549 261585 234583
rect 261585 234549 261619 234583
rect 261619 234549 261628 234583
rect 261576 234540 261628 234549
rect 246488 234472 246540 234524
rect 231216 231820 231268 231872
rect 231400 231820 231452 231872
rect 331772 231820 331824 231872
rect 335820 231820 335872 231872
rect 331864 231752 331916 231804
rect 335912 231752 335964 231804
rect 253020 230528 253072 230580
rect 253112 230528 253164 230580
rect 340144 230528 340196 230580
rect 107476 230460 107528 230512
rect 107660 230460 107712 230512
rect 232044 230503 232096 230512
rect 232044 230469 232053 230503
rect 232053 230469 232087 230503
rect 232087 230469 232096 230503
rect 232044 230460 232096 230469
rect 237840 230460 237892 230512
rect 237932 230460 237984 230512
rect 240508 230460 240560 230512
rect 240692 230460 240744 230512
rect 257068 230460 257120 230512
rect 257160 230460 257212 230512
rect 320916 230460 320968 230512
rect 321100 230460 321152 230512
rect 326252 230460 326304 230512
rect 326344 230460 326396 230512
rect 339960 230460 340012 230512
rect 330760 230052 330812 230104
rect 260196 229168 260248 229220
rect 260380 229168 260432 229220
rect 260380 229075 260432 229084
rect 260380 229041 260389 229075
rect 260389 229041 260423 229075
rect 260423 229041 260432 229075
rect 260380 229032 260432 229041
rect 340144 229032 340196 229084
rect 299020 227783 299072 227792
rect 299020 227749 299029 227783
rect 299029 227749 299063 227783
rect 299063 227749 299072 227783
rect 299020 227740 299072 227749
rect 300308 227715 300360 227724
rect 300308 227681 300317 227715
rect 300317 227681 300351 227715
rect 300351 227681 300360 227715
rect 300308 227672 300360 227681
rect 333060 227715 333112 227724
rect 333060 227681 333069 227715
rect 333069 227681 333103 227715
rect 333103 227681 333112 227715
rect 333060 227672 333112 227681
rect 299020 227647 299072 227656
rect 299020 227613 299029 227647
rect 299029 227613 299063 227647
rect 299063 227613 299072 227647
rect 299020 227604 299072 227613
rect 267188 227060 267240 227112
rect 268660 227060 268712 227112
rect 267188 226924 267240 226976
rect 268660 226924 268712 226976
rect 301780 226355 301832 226364
rect 301780 226321 301789 226355
rect 301789 226321 301823 226355
rect 301823 226321 301832 226355
rect 301780 226312 301832 226321
rect 232044 224995 232096 225004
rect 232044 224961 232053 224995
rect 232053 224961 232087 224995
rect 232087 224961 232096 224995
rect 232044 224952 232096 224961
rect 257068 224952 257120 225004
rect 344100 224952 344152 225004
rect 344284 224952 344336 225004
rect 257160 224884 257212 224936
rect 330760 224884 330812 224936
rect 330944 224884 330996 224936
rect 260380 224247 260432 224256
rect 260380 224213 260389 224247
rect 260389 224213 260423 224247
rect 260423 224213 260432 224247
rect 260380 224204 260432 224213
rect 322112 224204 322164 224256
rect 322296 224204 322348 224256
rect 2780 223048 2832 223100
rect 5172 223048 5224 223100
rect 232320 222232 232372 222284
rect 232596 222232 232648 222284
rect 100668 222164 100720 222216
rect 100852 222164 100904 222216
rect 232044 222207 232096 222216
rect 232044 222173 232053 222207
rect 232053 222173 232087 222207
rect 232087 222173 232096 222207
rect 232044 222164 232096 222173
rect 237932 222164 237984 222216
rect 238024 222164 238076 222216
rect 331772 222164 331824 222216
rect 331864 222164 331916 222216
rect 333244 222164 333296 222216
rect 333336 222164 333388 222216
rect 326344 220872 326396 220924
rect 253112 220804 253164 220856
rect 253296 220804 253348 220856
rect 293132 220804 293184 220856
rect 293316 220804 293368 220856
rect 320916 220804 320968 220856
rect 321100 220804 321152 220856
rect 326252 220804 326304 220856
rect 340052 220779 340104 220788
rect 340052 220745 340061 220779
rect 340061 220745 340095 220779
rect 340095 220745 340104 220779
rect 340052 220736 340104 220745
rect 260380 219419 260432 219428
rect 260380 219385 260389 219419
rect 260389 219385 260423 219419
rect 260423 219385 260432 219419
rect 260380 219376 260432 219385
rect 261576 219419 261628 219428
rect 261576 219385 261585 219419
rect 261585 219385 261619 219419
rect 261619 219385 261628 219419
rect 261576 219376 261628 219385
rect 265624 219376 265676 219428
rect 265808 219376 265860 219428
rect 319628 219419 319680 219428
rect 319628 219385 319637 219419
rect 319637 219385 319671 219419
rect 319671 219385 319680 219419
rect 319628 219376 319680 219385
rect 321100 219419 321152 219428
rect 321100 219385 321109 219419
rect 321109 219385 321143 219419
rect 321143 219385 321152 219419
rect 321100 219376 321152 219385
rect 322296 219308 322348 219360
rect 299020 218059 299072 218068
rect 299020 218025 299029 218059
rect 299029 218025 299063 218059
rect 299063 218025 299072 218059
rect 299020 218016 299072 218025
rect 300308 218059 300360 218068
rect 300308 218025 300317 218059
rect 300317 218025 300351 218059
rect 300351 218025 300360 218059
rect 300308 218016 300360 218025
rect 333152 218016 333204 218068
rect 335820 218016 335872 218068
rect 335912 218016 335964 218068
rect 333244 217948 333296 218000
rect 333336 217880 333388 217932
rect 246488 217404 246540 217456
rect 301780 216631 301832 216640
rect 301780 216597 301789 216631
rect 301789 216597 301823 216631
rect 301823 216597 301832 216631
rect 301780 216588 301832 216597
rect 334532 216588 334584 216640
rect 341708 215976 341760 216028
rect 341892 215976 341944 216028
rect 326252 215407 326304 215416
rect 326252 215373 326261 215407
rect 326261 215373 326295 215407
rect 326295 215373 326304 215407
rect 326252 215364 326304 215373
rect 261576 215271 261628 215280
rect 261576 215237 261585 215271
rect 261585 215237 261619 215271
rect 261619 215237 261628 215271
rect 261576 215228 261628 215237
rect 329012 215271 329064 215280
rect 329012 215237 329021 215271
rect 329021 215237 329055 215271
rect 329055 215237 329064 215271
rect 329012 215228 329064 215237
rect 330760 215228 330812 215280
rect 330944 215228 330996 215280
rect 232596 215092 232648 215144
rect 232780 215092 232832 215144
rect 260380 214523 260432 214532
rect 260380 214489 260389 214523
rect 260389 214489 260423 214523
rect 260423 214489 260432 214523
rect 260380 214480 260432 214489
rect 245016 212644 245068 212696
rect 231216 212508 231268 212560
rect 231400 212508 231452 212560
rect 245016 212440 245068 212492
rect 240692 211080 240744 211132
rect 240876 211080 240928 211132
rect 264336 211080 264388 211132
rect 264520 211080 264572 211132
rect 293132 211080 293184 211132
rect 293316 211080 293368 211132
rect 294604 211080 294656 211132
rect 294788 211080 294840 211132
rect 295892 211080 295944 211132
rect 296076 211080 296128 211132
rect 340052 211123 340104 211132
rect 340052 211089 340061 211123
rect 340061 211089 340095 211123
rect 340095 211089 340104 211123
rect 340052 211080 340104 211089
rect 246396 209831 246448 209840
rect 246396 209797 246405 209831
rect 246405 209797 246439 209831
rect 246439 209797 246448 209831
rect 246396 209788 246448 209797
rect 319628 209831 319680 209840
rect 319628 209797 319637 209831
rect 319637 209797 319671 209831
rect 319671 209797 319680 209831
rect 319628 209788 319680 209797
rect 321100 209831 321152 209840
rect 321100 209797 321109 209831
rect 321109 209797 321143 209831
rect 321143 209797 321152 209831
rect 321100 209788 321152 209797
rect 322112 209831 322164 209840
rect 322112 209797 322121 209831
rect 322121 209797 322155 209831
rect 322155 209797 322164 209831
rect 322112 209788 322164 209797
rect 335820 209763 335872 209772
rect 335820 209729 335829 209763
rect 335829 209729 335863 209763
rect 335863 209729 335872 209763
rect 335820 209720 335872 209729
rect 299020 208496 299072 208548
rect 331772 208428 331824 208480
rect 299020 208360 299072 208412
rect 331864 208360 331916 208412
rect 300308 208335 300360 208344
rect 300308 208301 300317 208335
rect 300317 208301 300351 208335
rect 300351 208301 300360 208335
rect 300308 208292 300360 208301
rect 267188 207748 267240 207800
rect 268660 207748 268712 207800
rect 267188 207612 267240 207664
rect 268660 207612 268712 207664
rect 301596 207000 301648 207052
rect 334624 207043 334676 207052
rect 334624 207009 334633 207043
rect 334633 207009 334667 207043
rect 334667 207009 334676 207043
rect 334624 207000 334676 207009
rect 246396 205640 246448 205692
rect 329104 205640 329156 205692
rect 344100 205640 344152 205692
rect 344284 205640 344336 205692
rect 262864 205572 262916 205624
rect 263048 205572 263100 205624
rect 330760 205572 330812 205624
rect 246488 205504 246540 205556
rect 340236 204892 340288 204944
rect 261576 203600 261628 203652
rect 261668 203600 261720 203652
rect 336096 203532 336148 203584
rect 244556 202920 244608 202972
rect 100668 202852 100720 202904
rect 100852 202852 100904 202904
rect 232320 202852 232372 202904
rect 232596 202852 232648 202904
rect 238024 202852 238076 202904
rect 238116 202852 238168 202904
rect 244464 202895 244516 202904
rect 244464 202861 244473 202895
rect 244473 202861 244507 202895
rect 244507 202861 244516 202895
rect 244464 202852 244516 202861
rect 257160 202920 257212 202972
rect 253020 202852 253072 202904
rect 253112 202852 253164 202904
rect 257068 202852 257120 202904
rect 258724 202852 258776 202904
rect 258816 202852 258868 202904
rect 260288 202852 260340 202904
rect 260380 202852 260432 202904
rect 244556 202784 244608 202836
rect 244464 201535 244516 201544
rect 244464 201501 244473 201535
rect 244473 201501 244507 201535
rect 244507 201501 244516 201535
rect 244464 201492 244516 201501
rect 107476 201424 107528 201476
rect 107660 201424 107712 201476
rect 264336 201424 264388 201476
rect 264520 201424 264572 201476
rect 293132 201424 293184 201476
rect 293316 201424 293368 201476
rect 345388 201424 345440 201476
rect 345572 201424 345624 201476
rect 326252 200175 326304 200184
rect 326252 200141 326261 200175
rect 326261 200141 326295 200175
rect 326295 200141 326304 200175
rect 326252 200132 326304 200141
rect 319628 200107 319680 200116
rect 319628 200073 319637 200107
rect 319637 200073 319671 200107
rect 319671 200073 319680 200107
rect 319628 200064 319680 200073
rect 321100 200107 321152 200116
rect 321100 200073 321109 200107
rect 321109 200073 321143 200107
rect 321143 200073 321152 200107
rect 321100 200064 321152 200073
rect 322296 200064 322348 200116
rect 300308 198747 300360 198756
rect 300308 198713 300317 198747
rect 300317 198713 300351 198747
rect 300351 198713 300360 198747
rect 300308 198704 300360 198713
rect 299020 198679 299072 198688
rect 299020 198645 299029 198679
rect 299029 198645 299063 198679
rect 299063 198645 299072 198679
rect 299020 198636 299072 198645
rect 301780 197276 301832 197328
rect 329104 197276 329156 197328
rect 331864 197276 331916 197328
rect 332048 197276 332100 197328
rect 334624 197319 334676 197328
rect 334624 197285 334633 197319
rect 334633 197285 334667 197319
rect 334667 197285 334676 197319
rect 334624 197276 334676 197285
rect 326252 196052 326304 196104
rect 232780 195984 232832 196036
rect 232688 195916 232740 195968
rect 326252 195916 326304 195968
rect 341524 195916 341576 195968
rect 341708 195916 341760 195968
rect 245016 195236 245068 195288
rect 2780 194284 2832 194336
rect 5080 194284 5132 194336
rect 231216 193196 231268 193248
rect 231400 193196 231452 193248
rect 232320 193196 232372 193248
rect 232412 193196 232464 193248
rect 246396 193196 246448 193248
rect 246580 193196 246632 193248
rect 333060 193196 333112 193248
rect 333152 193196 333204 193248
rect 253020 191836 253072 191888
rect 253112 191836 253164 191888
rect 258816 191836 258868 191888
rect 258908 191836 258960 191888
rect 232136 191768 232188 191820
rect 232412 191768 232464 191820
rect 240692 191768 240744 191820
rect 260196 191811 260248 191820
rect 260196 191777 260205 191811
rect 260205 191777 260239 191811
rect 260239 191777 260248 191811
rect 260196 191768 260248 191777
rect 264336 191768 264388 191820
rect 264520 191768 264572 191820
rect 265624 191768 265676 191820
rect 265808 191768 265860 191820
rect 293132 191768 293184 191820
rect 293316 191768 293368 191820
rect 294604 191768 294656 191820
rect 294788 191768 294840 191820
rect 295892 191768 295944 191820
rect 296076 191768 296128 191820
rect 333060 191768 333112 191820
rect 333152 191768 333204 191820
rect 240876 191700 240928 191752
rect 319628 190519 319680 190528
rect 319628 190485 319637 190519
rect 319637 190485 319671 190519
rect 319671 190485 319680 190519
rect 319628 190476 319680 190485
rect 321100 190519 321152 190528
rect 321100 190485 321109 190519
rect 321109 190485 321143 190519
rect 321143 190485 321152 190519
rect 321100 190476 321152 190485
rect 322204 190519 322256 190528
rect 322204 190485 322213 190519
rect 322213 190485 322247 190519
rect 322247 190485 322256 190519
rect 322204 190476 322256 190485
rect 261484 190451 261536 190460
rect 261484 190417 261493 190451
rect 261493 190417 261527 190451
rect 261527 190417 261536 190451
rect 261484 190408 261536 190417
rect 263048 190451 263100 190460
rect 263048 190417 263057 190451
rect 263057 190417 263091 190451
rect 263091 190417 263100 190451
rect 263048 190408 263100 190417
rect 333244 190408 333296 190460
rect 333336 190408 333388 190460
rect 335820 190451 335872 190460
rect 335820 190417 335829 190451
rect 335829 190417 335863 190451
rect 335863 190417 335872 190451
rect 335820 190408 335872 190417
rect 244188 189456 244240 189508
rect 299020 189091 299072 189100
rect 299020 189057 299029 189091
rect 299029 189057 299063 189091
rect 299063 189057 299072 189091
rect 299020 189048 299072 189057
rect 300308 189023 300360 189032
rect 300308 188989 300317 189023
rect 300317 188989 300351 189023
rect 300351 188989 300360 189023
rect 300308 188980 300360 188989
rect 301780 187731 301832 187740
rect 301780 187697 301789 187731
rect 301789 187697 301823 187731
rect 301823 187697 301832 187731
rect 301780 187688 301832 187697
rect 329012 187731 329064 187740
rect 329012 187697 329021 187731
rect 329021 187697 329055 187731
rect 329055 187697 329064 187731
rect 329012 187688 329064 187697
rect 330576 187731 330628 187740
rect 330576 187697 330585 187731
rect 330585 187697 330619 187731
rect 330619 187697 330628 187731
rect 330576 187688 330628 187697
rect 334624 187731 334676 187740
rect 334624 187697 334633 187731
rect 334633 187697 334667 187731
rect 334667 187697 334676 187731
rect 334624 187688 334676 187697
rect 257160 186396 257212 186448
rect 258908 186328 258960 186380
rect 257068 186260 257120 186312
rect 258908 186192 258960 186244
rect 333152 183923 333204 183932
rect 333152 183889 333161 183923
rect 333161 183889 333195 183923
rect 333195 183889 333204 183923
rect 333152 183880 333204 183889
rect 345388 183608 345440 183660
rect 100668 183540 100720 183592
rect 100852 183540 100904 183592
rect 238024 183540 238076 183592
rect 238116 183540 238168 183592
rect 245016 183540 245068 183592
rect 341616 183540 341668 183592
rect 341708 183540 341760 183592
rect 345296 183540 345348 183592
rect 260288 183472 260340 183524
rect 107476 182112 107528 182164
rect 107660 182112 107712 182164
rect 232044 182112 232096 182164
rect 232320 182155 232372 182164
rect 232320 182121 232329 182155
rect 232329 182121 232363 182155
rect 232363 182121 232372 182155
rect 232320 182112 232372 182121
rect 260288 182155 260340 182164
rect 260288 182121 260297 182155
rect 260297 182121 260331 182155
rect 260331 182121 260340 182155
rect 260288 182112 260340 182121
rect 261484 182155 261536 182164
rect 261484 182121 261493 182155
rect 261493 182121 261527 182155
rect 261527 182121 261536 182155
rect 261484 182112 261536 182121
rect 293132 182112 293184 182164
rect 293316 182112 293368 182164
rect 231952 182044 232004 182096
rect 333152 182087 333204 182096
rect 333152 182053 333161 182087
rect 333161 182053 333195 182087
rect 333195 182053 333204 182087
rect 333152 182044 333204 182053
rect 263048 180863 263100 180872
rect 263048 180829 263057 180863
rect 263057 180829 263091 180863
rect 263091 180829 263100 180863
rect 263048 180820 263100 180829
rect 334624 180820 334676 180872
rect 335820 180863 335872 180872
rect 335820 180829 335829 180863
rect 335829 180829 335863 180863
rect 335863 180829 335872 180863
rect 335820 180820 335872 180829
rect 264520 180795 264572 180804
rect 264520 180761 264529 180795
rect 264529 180761 264563 180795
rect 264563 180761 264572 180795
rect 264520 180752 264572 180761
rect 265808 180795 265860 180804
rect 265808 180761 265817 180795
rect 265817 180761 265851 180795
rect 265851 180761 265860 180795
rect 265808 180752 265860 180761
rect 293132 180795 293184 180804
rect 293132 180761 293141 180795
rect 293141 180761 293175 180795
rect 293175 180761 293184 180795
rect 293132 180752 293184 180761
rect 319628 180795 319680 180804
rect 319628 180761 319637 180795
rect 319637 180761 319671 180795
rect 319671 180761 319680 180795
rect 319628 180752 319680 180761
rect 321100 180795 321152 180804
rect 321100 180761 321109 180795
rect 321109 180761 321143 180795
rect 321143 180761 321152 180795
rect 321100 180752 321152 180761
rect 2780 179664 2832 179716
rect 4988 179664 5040 179716
rect 301780 179596 301832 179648
rect 301780 179460 301832 179512
rect 334532 179503 334584 179512
rect 334532 179469 334541 179503
rect 334541 179469 334575 179503
rect 334575 179469 334584 179503
rect 334532 179460 334584 179469
rect 298928 179392 298980 179444
rect 299020 179392 299072 179444
rect 300308 179435 300360 179444
rect 300308 179401 300317 179435
rect 300317 179401 300351 179435
rect 300351 179401 300360 179435
rect 300308 179392 300360 179401
rect 329012 179324 329064 179376
rect 329104 179324 329156 179376
rect 334532 179367 334584 179376
rect 334532 179333 334541 179367
rect 334541 179333 334575 179367
rect 334575 179333 334584 179367
rect 334532 179324 334584 179333
rect 340052 178780 340104 178832
rect 340144 178712 340196 178764
rect 331864 178032 331916 178084
rect 332048 178032 332100 178084
rect 301780 178007 301832 178016
rect 301780 177973 301789 178007
rect 301789 177973 301823 178007
rect 301823 177973 301832 178007
rect 301780 177964 301832 177973
rect 232688 176604 232740 176656
rect 232688 176468 232740 176520
rect 231216 173884 231268 173936
rect 231400 173884 231452 173936
rect 244464 173884 244516 173936
rect 244924 173884 244976 173936
rect 245108 173884 245160 173936
rect 245844 173884 245896 173936
rect 246028 173884 246080 173936
rect 246396 173884 246448 173936
rect 246580 173884 246632 173936
rect 333244 173884 333296 173936
rect 335820 173884 335872 173936
rect 345296 173884 345348 173936
rect 345388 173884 345440 173936
rect 260288 173859 260340 173868
rect 260288 173825 260297 173859
rect 260297 173825 260331 173859
rect 260331 173825 260340 173859
rect 260288 173816 260340 173825
rect 333336 173748 333388 173800
rect 335912 173748 335964 173800
rect 232412 172524 232464 172576
rect 252928 172524 252980 172576
rect 253020 172524 253072 172576
rect 256976 172524 257028 172576
rect 257068 172524 257120 172576
rect 258816 172524 258868 172576
rect 258908 172524 258960 172576
rect 240692 172456 240744 172508
rect 240876 172456 240928 172508
rect 294788 171232 294840 171284
rect 296076 171232 296128 171284
rect 322296 171164 322348 171216
rect 264520 171139 264572 171148
rect 264520 171105 264529 171139
rect 264529 171105 264563 171139
rect 264563 171105 264572 171139
rect 264520 171096 264572 171105
rect 265808 171139 265860 171148
rect 265808 171105 265817 171139
rect 265817 171105 265851 171139
rect 265851 171105 265860 171139
rect 265808 171096 265860 171105
rect 293316 171096 293368 171148
rect 294788 171096 294840 171148
rect 296076 171096 296128 171148
rect 319628 171139 319680 171148
rect 319628 171105 319637 171139
rect 319637 171105 319671 171139
rect 319671 171105 319680 171139
rect 319628 171096 319680 171105
rect 321100 171139 321152 171148
rect 321100 171105 321109 171139
rect 321109 171105 321143 171139
rect 321143 171105 321152 171139
rect 321100 171096 321152 171105
rect 322388 171096 322440 171148
rect 334532 171071 334584 171080
rect 334532 171037 334541 171071
rect 334541 171037 334575 171071
rect 334575 171037 334584 171071
rect 334532 171028 334584 171037
rect 331864 169804 331916 169856
rect 299020 169711 299072 169720
rect 299020 169677 299029 169711
rect 299029 169677 299063 169711
rect 299063 169677 299072 169711
rect 299020 169668 299072 169677
rect 300308 169711 300360 169720
rect 300308 169677 300317 169711
rect 300317 169677 300351 169711
rect 300351 169677 300360 169711
rect 300308 169668 300360 169677
rect 326344 169711 326396 169720
rect 326344 169677 326353 169711
rect 326353 169677 326387 169711
rect 326387 169677 326396 169711
rect 326344 169668 326396 169677
rect 340144 169056 340196 169108
rect 340328 169056 340380 169108
rect 301780 168419 301832 168428
rect 301780 168385 301789 168419
rect 301789 168385 301823 168419
rect 301823 168385 301832 168419
rect 301780 168376 301832 168385
rect 331772 168419 331824 168428
rect 331772 168385 331781 168419
rect 331781 168385 331815 168419
rect 331815 168385 331824 168419
rect 331772 168376 331824 168385
rect 231952 167628 232004 167680
rect 232136 167628 232188 167680
rect 322388 167084 322440 167136
rect 232412 167016 232464 167068
rect 232320 166948 232372 167000
rect 322296 166880 322348 166932
rect 335912 166268 335964 166320
rect 336096 166268 336148 166320
rect 261668 164296 261720 164348
rect 252928 164228 252980 164280
rect 253020 164228 253072 164280
rect 256976 164228 257028 164280
rect 257068 164228 257120 164280
rect 261576 164228 261628 164280
rect 244188 164160 244240 164212
rect 244372 164160 244424 164212
rect 340052 164160 340104 164212
rect 340144 164160 340196 164212
rect 345388 164160 345440 164212
rect 345572 164160 345624 164212
rect 107476 162843 107528 162852
rect 107476 162809 107485 162843
rect 107485 162809 107519 162843
rect 107519 162809 107528 162843
rect 107476 162800 107528 162809
rect 232044 162800 232096 162852
rect 232136 162800 232188 162852
rect 232320 162800 232372 162852
rect 232596 162800 232648 162852
rect 261576 162800 261628 162852
rect 261668 162800 261720 162852
rect 329012 161440 329064 161492
rect 329104 161440 329156 161492
rect 232596 161415 232648 161424
rect 232596 161381 232605 161415
rect 232605 161381 232639 161415
rect 232639 161381 232648 161415
rect 232596 161372 232648 161381
rect 253020 161415 253072 161424
rect 253020 161381 253029 161415
rect 253029 161381 253063 161415
rect 253063 161381 253072 161415
rect 253020 161372 253072 161381
rect 257068 161415 257120 161424
rect 257068 161381 257077 161415
rect 257077 161381 257111 161415
rect 257111 161381 257120 161415
rect 257068 161372 257120 161381
rect 293316 161415 293368 161424
rect 293316 161381 293325 161415
rect 293325 161381 293359 161415
rect 293359 161381 293368 161415
rect 293316 161372 293368 161381
rect 319628 161415 319680 161424
rect 319628 161381 319637 161415
rect 319637 161381 319671 161415
rect 319671 161381 319680 161415
rect 319628 161372 319680 161381
rect 321100 161415 321152 161424
rect 321100 161381 321109 161415
rect 321109 161381 321143 161415
rect 321143 161381 321152 161415
rect 321100 161372 321152 161381
rect 326436 161304 326488 161356
rect 301872 160352 301924 160404
rect 299020 160123 299072 160132
rect 299020 160089 299029 160123
rect 299029 160089 299063 160123
rect 299063 160089 299072 160123
rect 299020 160080 299072 160089
rect 300308 160123 300360 160132
rect 300308 160089 300317 160123
rect 300317 160089 300351 160123
rect 300351 160089 300360 160123
rect 300308 160080 300360 160089
rect 301780 160080 301832 160132
rect 301872 160080 301924 160132
rect 330484 160080 330536 160132
rect 330576 160080 330628 160132
rect 260380 160012 260432 160064
rect 260288 159944 260340 159996
rect 301780 159944 301832 159996
rect 260288 158695 260340 158704
rect 260288 158661 260297 158695
rect 260297 158661 260331 158695
rect 260331 158661 260340 158695
rect 260288 158652 260340 158661
rect 258816 157428 258868 157480
rect 231216 157292 231268 157344
rect 258816 157292 258868 157344
rect 231216 157156 231268 157208
rect 100668 154504 100720 154556
rect 100852 154504 100904 154556
rect 231216 154504 231268 154556
rect 231400 154504 231452 154556
rect 107476 153255 107528 153264
rect 107476 153221 107485 153255
rect 107485 153221 107519 153255
rect 107519 153221 107528 153255
rect 107476 153212 107528 153221
rect 257252 153212 257304 153264
rect 232136 153144 232188 153196
rect 232596 153187 232648 153196
rect 232596 153153 232605 153187
rect 232605 153153 232639 153187
rect 232639 153153 232648 153187
rect 232596 153144 232648 153153
rect 240692 153144 240744 153196
rect 240876 153144 240928 153196
rect 257252 153076 257304 153128
rect 294788 151920 294840 151972
rect 296076 151920 296128 151972
rect 253020 151827 253072 151836
rect 253020 151793 253029 151827
rect 253029 151793 253063 151827
rect 253063 151793 253072 151827
rect 253020 151784 253072 151793
rect 257344 151784 257396 151836
rect 293316 151827 293368 151836
rect 293316 151793 293325 151827
rect 293325 151793 293359 151827
rect 293359 151793 293368 151827
rect 293316 151784 293368 151793
rect 294788 151784 294840 151836
rect 296076 151784 296128 151836
rect 319628 151827 319680 151836
rect 319628 151793 319637 151827
rect 319637 151793 319671 151827
rect 319671 151793 319680 151827
rect 319628 151784 319680 151793
rect 321100 151827 321152 151836
rect 321100 151793 321109 151827
rect 321109 151793 321143 151827
rect 321143 151793 321152 151827
rect 321100 151784 321152 151793
rect 333244 151784 333296 151836
rect 333336 151784 333388 151836
rect 264520 151759 264572 151768
rect 264520 151725 264529 151759
rect 264529 151725 264563 151759
rect 264563 151725 264572 151759
rect 264520 151716 264572 151725
rect 322296 151716 322348 151768
rect 322388 151716 322440 151768
rect 331772 151759 331824 151768
rect 331772 151725 331781 151759
rect 331781 151725 331815 151759
rect 331815 151725 331824 151759
rect 331772 151716 331824 151725
rect 334532 151759 334584 151768
rect 334532 151725 334541 151759
rect 334541 151725 334575 151759
rect 334575 151725 334584 151759
rect 334532 151716 334584 151725
rect 253020 151691 253072 151700
rect 253020 151657 253029 151691
rect 253029 151657 253063 151691
rect 253063 151657 253072 151691
rect 253020 151648 253072 151657
rect 2780 151308 2832 151360
rect 4896 151308 4948 151360
rect 296076 150399 296128 150408
rect 296076 150365 296085 150399
rect 296085 150365 296119 150399
rect 296119 150365 296128 150399
rect 296076 150356 296128 150365
rect 330484 150399 330536 150408
rect 330484 150365 330493 150399
rect 330493 150365 330527 150399
rect 330527 150365 330536 150399
rect 330484 150356 330536 150365
rect 301780 150220 301832 150272
rect 260288 149107 260340 149116
rect 260288 149073 260297 149107
rect 260297 149073 260331 149107
rect 260331 149073 260340 149107
rect 260288 149064 260340 149073
rect 244464 147704 244516 147756
rect 244924 147704 244976 147756
rect 301504 147679 301556 147688
rect 301504 147645 301513 147679
rect 301513 147645 301547 147679
rect 301547 147645 301556 147679
rect 301504 147636 301556 147645
rect 344100 147636 344152 147688
rect 344284 147636 344336 147688
rect 244372 147568 244424 147620
rect 244924 147568 244976 147620
rect 345296 144916 345348 144968
rect 345388 144916 345440 144968
rect 232044 143599 232096 143608
rect 232044 143565 232053 143599
rect 232053 143565 232087 143599
rect 232087 143565 232096 143599
rect 232044 143556 232096 143565
rect 246396 143599 246448 143608
rect 246396 143565 246405 143599
rect 246405 143565 246439 143599
rect 246439 143565 246448 143599
rect 246396 143556 246448 143565
rect 320916 143556 320968 143608
rect 321100 143556 321152 143608
rect 107476 143531 107528 143540
rect 107476 143497 107485 143531
rect 107485 143497 107519 143531
rect 107519 143497 107528 143531
rect 107476 143488 107528 143497
rect 240692 143531 240744 143540
rect 240692 143497 240701 143531
rect 240701 143497 240735 143531
rect 240735 143497 240744 143531
rect 240692 143488 240744 143497
rect 244372 143488 244424 143540
rect 244464 143488 244516 143540
rect 246028 143531 246080 143540
rect 246028 143497 246037 143531
rect 246037 143497 246071 143531
rect 246071 143497 246080 143531
rect 246028 143488 246080 143497
rect 254676 143488 254728 143540
rect 254860 143488 254912 143540
rect 258816 143531 258868 143540
rect 258816 143497 258825 143531
rect 258825 143497 258859 143531
rect 258859 143497 258868 143531
rect 258816 143488 258868 143497
rect 314292 143488 314344 143540
rect 314384 143531 314436 143540
rect 314384 143497 314393 143531
rect 314393 143497 314427 143531
rect 314427 143497 314436 143531
rect 314384 143488 314436 143497
rect 314200 143420 314252 143472
rect 314292 143352 314344 143404
rect 314200 143284 314252 143336
rect 253204 142196 253256 142248
rect 246396 142171 246448 142180
rect 246396 142137 246405 142171
rect 246405 142137 246439 142171
rect 246439 142137 246448 142171
rect 246396 142128 246448 142137
rect 256976 142128 257028 142180
rect 257344 142128 257396 142180
rect 260288 142128 260340 142180
rect 264520 142171 264572 142180
rect 264520 142137 264529 142171
rect 264529 142137 264563 142171
rect 264563 142137 264572 142171
rect 264520 142128 264572 142137
rect 294696 142128 294748 142180
rect 294788 142128 294840 142180
rect 326160 142128 326212 142180
rect 326344 142128 326396 142180
rect 331772 142171 331824 142180
rect 331772 142137 331781 142171
rect 331781 142137 331815 142171
rect 331815 142137 331824 142171
rect 331772 142128 331824 142137
rect 334532 142171 334584 142180
rect 334532 142137 334541 142171
rect 334541 142137 334575 142171
rect 334575 142137 334584 142171
rect 334532 142128 334584 142137
rect 232044 142103 232096 142112
rect 232044 142069 232053 142103
rect 232053 142069 232087 142103
rect 232087 142069 232096 142103
rect 232044 142060 232096 142069
rect 293316 142103 293368 142112
rect 293316 142069 293325 142103
rect 293325 142069 293359 142103
rect 293359 142069 293368 142103
rect 293316 142060 293368 142069
rect 319628 142103 319680 142112
rect 319628 142069 319637 142103
rect 319637 142069 319671 142103
rect 319671 142069 319680 142103
rect 319628 142060 319680 142069
rect 322296 142060 322348 142112
rect 246396 141992 246448 142044
rect 260288 141992 260340 142044
rect 322296 141924 322348 141976
rect 301872 141083 301924 141092
rect 301872 141049 301881 141083
rect 301881 141049 301915 141083
rect 301915 141049 301924 141083
rect 301872 141040 301924 141049
rect 296168 140768 296220 140820
rect 330392 140768 330444 140820
rect 244924 140743 244976 140752
rect 244924 140709 244933 140743
rect 244933 140709 244967 140743
rect 244967 140709 244976 140743
rect 244924 140700 244976 140709
rect 253204 140743 253256 140752
rect 253204 140709 253213 140743
rect 253213 140709 253247 140743
rect 253247 140709 253256 140743
rect 253204 140700 253256 140709
rect 299020 140743 299072 140752
rect 299020 140709 299029 140743
rect 299029 140709 299063 140743
rect 299063 140709 299072 140743
rect 299020 140700 299072 140709
rect 300308 140743 300360 140752
rect 300308 140709 300317 140743
rect 300317 140709 300351 140743
rect 300351 140709 300360 140743
rect 300308 140700 300360 140709
rect 301504 140700 301556 140752
rect 301780 140700 301832 140752
rect 329012 140743 329064 140752
rect 329012 140709 329021 140743
rect 329021 140709 329055 140743
rect 329055 140709 329064 140743
rect 329012 140700 329064 140709
rect 331772 140743 331824 140752
rect 331772 140709 331781 140743
rect 331781 140709 331815 140743
rect 331815 140709 331824 140743
rect 331772 140700 331824 140709
rect 335820 140700 335872 140752
rect 301872 140675 301924 140684
rect 301872 140641 301881 140675
rect 301881 140641 301915 140675
rect 301915 140641 301924 140675
rect 301872 140632 301924 140641
rect 232412 139340 232464 139392
rect 232596 139340 232648 139392
rect 260196 139383 260248 139392
rect 260196 139349 260205 139383
rect 260205 139349 260239 139383
rect 260239 139349 260248 139383
rect 260196 139340 260248 139349
rect 258908 138592 258960 138644
rect 314384 138499 314436 138508
rect 314384 138465 314393 138499
rect 314393 138465 314427 138499
rect 314427 138465 314436 138499
rect 314384 138456 314436 138465
rect 232596 138048 232648 138100
rect 232688 138048 232740 138100
rect 231216 138023 231268 138032
rect 231216 137989 231225 138023
rect 231225 137989 231259 138023
rect 231259 137989 231268 138023
rect 231216 137980 231268 137989
rect 232412 136552 232464 136604
rect 2780 136348 2832 136400
rect 4804 136348 4856 136400
rect 231216 135371 231268 135380
rect 231216 135337 231225 135371
rect 231225 135337 231259 135371
rect 231259 135337 231268 135371
rect 231216 135328 231268 135337
rect 340144 135260 340196 135312
rect 345296 135260 345348 135312
rect 345388 135260 345440 135312
rect 100668 135192 100720 135244
rect 100852 135192 100904 135244
rect 231216 135192 231268 135244
rect 231400 135192 231452 135244
rect 340052 135192 340104 135244
rect 301780 134555 301832 134564
rect 301780 134521 301789 134555
rect 301789 134521 301823 134555
rect 301823 134521 301832 134555
rect 301780 134512 301832 134521
rect 107476 133943 107528 133952
rect 107476 133909 107485 133943
rect 107485 133909 107519 133943
rect 107519 133909 107528 133943
rect 107476 133900 107528 133909
rect 240692 133943 240744 133952
rect 240692 133909 240701 133943
rect 240701 133909 240735 133943
rect 240735 133909 240744 133943
rect 240692 133900 240744 133909
rect 340052 133875 340104 133884
rect 340052 133841 340061 133875
rect 340061 133841 340095 133875
rect 340095 133841 340104 133875
rect 340052 133832 340104 133841
rect 345388 133832 345440 133884
rect 345572 133832 345624 133884
rect 245844 133288 245896 133340
rect 232136 132472 232188 132524
rect 293316 132515 293368 132524
rect 293316 132481 293325 132515
rect 293325 132481 293359 132515
rect 293359 132481 293368 132515
rect 293316 132472 293368 132481
rect 294788 132472 294840 132524
rect 294880 132472 294932 132524
rect 319628 132515 319680 132524
rect 319628 132481 319637 132515
rect 319637 132481 319671 132515
rect 319671 132481 319680 132515
rect 319628 132472 319680 132481
rect 321008 132472 321060 132524
rect 321100 132472 321152 132524
rect 326160 132472 326212 132524
rect 326252 132472 326304 132524
rect 330392 132472 330444 132524
rect 330484 132472 330536 132524
rect 261484 131180 261536 131232
rect 261576 131180 261628 131232
rect 245108 131112 245160 131164
rect 253204 131155 253256 131164
rect 253204 131121 253213 131155
rect 253213 131121 253247 131155
rect 253247 131121 253256 131155
rect 253204 131112 253256 131121
rect 329196 131112 329248 131164
rect 331772 131155 331824 131164
rect 331772 131121 331781 131155
rect 331781 131121 331815 131155
rect 331815 131121 331824 131155
rect 331772 131112 331824 131121
rect 335912 131155 335964 131164
rect 335912 131121 335921 131155
rect 335921 131121 335955 131155
rect 335955 131121 335964 131155
rect 335912 131112 335964 131121
rect 261484 131087 261536 131096
rect 261484 131053 261493 131087
rect 261493 131053 261527 131087
rect 261527 131053 261536 131087
rect 261484 131044 261536 131053
rect 334532 131044 334584 131096
rect 300308 130747 300360 130756
rect 300308 130713 300317 130747
rect 300317 130713 300351 130747
rect 300351 130713 300360 130747
rect 300308 130704 300360 130713
rect 299020 129863 299072 129872
rect 299020 129829 299029 129863
rect 299029 129829 299063 129863
rect 299063 129829 299072 129863
rect 299020 129820 299072 129829
rect 260288 129752 260340 129804
rect 299020 129727 299072 129736
rect 299020 129693 299029 129727
rect 299029 129693 299063 129727
rect 299063 129693 299072 129727
rect 299020 129684 299072 129693
rect 344100 128324 344152 128376
rect 344284 128324 344336 128376
rect 232872 127032 232924 127084
rect 232688 126964 232740 127016
rect 258816 125604 258868 125656
rect 258908 125604 258960 125656
rect 246396 124219 246448 124228
rect 246396 124185 246405 124219
rect 246405 124185 246439 124219
rect 246439 124185 246448 124219
rect 246396 124176 246448 124185
rect 326252 124176 326304 124228
rect 326344 124176 326396 124228
rect 329104 124176 329156 124228
rect 329196 124176 329248 124228
rect 340144 124176 340196 124228
rect 107476 124151 107528 124160
rect 107476 124117 107485 124151
rect 107485 124117 107519 124151
rect 107519 124117 107528 124151
rect 107476 124108 107528 124117
rect 317144 124151 317196 124160
rect 317144 124117 317153 124151
rect 317153 124117 317187 124151
rect 317187 124117 317196 124151
rect 317144 124108 317196 124117
rect 317328 124151 317380 124160
rect 317328 124117 317337 124151
rect 317337 124117 317371 124151
rect 317371 124117 317380 124151
rect 317328 124108 317380 124117
rect 345296 124108 345348 124160
rect 577504 124108 577556 124160
rect 579620 124108 579672 124160
rect 314384 124040 314436 124092
rect 345388 124040 345440 124092
rect 314384 123904 314436 123956
rect 321100 122884 321152 122936
rect 294696 122816 294748 122868
rect 294788 122816 294840 122868
rect 320916 122816 320968 122868
rect 244372 122791 244424 122800
rect 244372 122757 244381 122791
rect 244381 122757 244415 122791
rect 244415 122757 244424 122791
rect 244372 122748 244424 122757
rect 253020 122748 253072 122800
rect 254768 122748 254820 122800
rect 257160 122791 257212 122800
rect 257160 122757 257169 122791
rect 257169 122757 257203 122791
rect 257203 122757 257212 122791
rect 257160 122748 257212 122757
rect 264520 122748 264572 122800
rect 265808 122791 265860 122800
rect 265808 122757 265817 122791
rect 265817 122757 265851 122791
rect 265851 122757 265860 122791
rect 265808 122748 265860 122757
rect 319628 122748 319680 122800
rect 261484 122723 261536 122732
rect 261484 122689 261493 122723
rect 261493 122689 261527 122723
rect 261527 122689 261536 122723
rect 261484 122680 261536 122689
rect 322296 122884 322348 122936
rect 335728 122884 335780 122936
rect 335912 122884 335964 122936
rect 335728 122748 335780 122800
rect 335820 122748 335872 122800
rect 322388 122680 322440 122732
rect 301780 121499 301832 121508
rect 301780 121465 301789 121499
rect 301789 121465 301823 121499
rect 301823 121465 301832 121499
rect 301780 121456 301832 121465
rect 334532 121456 334584 121508
rect 245108 121388 245160 121440
rect 261484 121388 261536 121440
rect 331772 121431 331824 121440
rect 331772 121397 331781 121431
rect 331781 121397 331815 121431
rect 331815 121397 331824 121431
rect 331772 121388 331824 121397
rect 299020 120207 299072 120216
rect 299020 120173 299029 120207
rect 299029 120173 299063 120207
rect 299063 120173 299072 120207
rect 299020 120164 299072 120173
rect 299020 120028 299072 120080
rect 300308 120028 300360 120080
rect 301780 120028 301832 120080
rect 231216 118711 231268 118720
rect 231216 118677 231225 118711
rect 231225 118677 231259 118711
rect 231259 118677 231268 118711
rect 231216 118668 231268 118677
rect 232412 118711 232464 118720
rect 232412 118677 232421 118711
rect 232421 118677 232455 118711
rect 232455 118677 232464 118711
rect 232412 118668 232464 118677
rect 232596 118668 232648 118720
rect 232688 118668 232740 118720
rect 263048 118031 263100 118040
rect 263048 117997 263057 118031
rect 263057 117997 263091 118031
rect 263091 117997 263100 118031
rect 263048 117988 263100 117997
rect 317144 117555 317196 117564
rect 317144 117521 317153 117555
rect 317153 117521 317187 117555
rect 317187 117521 317196 117555
rect 317144 117512 317196 117521
rect 232688 117240 232740 117292
rect 232872 117172 232924 117224
rect 231216 116059 231268 116068
rect 231216 116025 231225 116059
rect 231225 116025 231259 116059
rect 231259 116025 231268 116059
rect 231216 116016 231268 116025
rect 100668 115923 100720 115932
rect 100668 115889 100677 115923
rect 100677 115889 100711 115923
rect 100711 115889 100720 115923
rect 100668 115880 100720 115889
rect 231216 115923 231268 115932
rect 231216 115889 231225 115923
rect 231225 115889 231259 115923
rect 231259 115889 231268 115923
rect 231216 115880 231268 115889
rect 258908 115923 258960 115932
rect 258908 115889 258917 115923
rect 258917 115889 258951 115923
rect 258951 115889 258960 115923
rect 258908 115880 258960 115889
rect 260380 115923 260432 115932
rect 260380 115889 260389 115923
rect 260389 115889 260423 115923
rect 260423 115889 260432 115923
rect 260380 115880 260432 115889
rect 317328 115583 317380 115592
rect 317328 115549 317337 115583
rect 317337 115549 317371 115583
rect 317371 115549 317380 115583
rect 317328 115540 317380 115549
rect 340144 115472 340196 115524
rect 107476 114563 107528 114572
rect 107476 114529 107485 114563
rect 107485 114529 107519 114563
rect 107519 114529 107528 114563
rect 107476 114520 107528 114529
rect 329012 114520 329064 114572
rect 329104 114520 329156 114572
rect 316960 114495 317012 114504
rect 316960 114461 316969 114495
rect 316969 114461 317003 114495
rect 317003 114461 317012 114495
rect 316960 114452 317012 114461
rect 317144 114495 317196 114504
rect 317144 114461 317153 114495
rect 317153 114461 317187 114495
rect 317187 114461 317196 114495
rect 317144 114452 317196 114461
rect 317328 114495 317380 114504
rect 317328 114461 317337 114495
rect 317337 114461 317371 114495
rect 317371 114461 317380 114495
rect 317328 114452 317380 114461
rect 326160 114452 326212 114504
rect 326344 114452 326396 114504
rect 317236 114427 317288 114436
rect 317236 114393 317245 114427
rect 317245 114393 317279 114427
rect 317279 114393 317288 114427
rect 317236 114384 317288 114393
rect 244464 113160 244516 113212
rect 257160 113203 257212 113212
rect 257160 113169 257169 113203
rect 257169 113169 257203 113203
rect 257203 113169 257212 113203
rect 257160 113160 257212 113169
rect 264520 113160 264572 113212
rect 265808 113203 265860 113212
rect 265808 113169 265817 113203
rect 265817 113169 265851 113203
rect 265851 113169 265860 113203
rect 265808 113160 265860 113169
rect 319628 113203 319680 113212
rect 319628 113169 319637 113203
rect 319637 113169 319671 113203
rect 319671 113169 319680 113203
rect 319628 113160 319680 113169
rect 245108 113092 245160 113144
rect 294788 113135 294840 113144
rect 294788 113101 294797 113135
rect 294797 113101 294831 113135
rect 294831 113101 294840 113135
rect 294788 113092 294840 113101
rect 326160 113135 326212 113144
rect 326160 113101 326169 113135
rect 326169 113101 326203 113135
rect 326203 113101 326212 113135
rect 326160 113092 326212 113101
rect 335820 113135 335872 113144
rect 335820 113101 335829 113135
rect 335829 113101 335863 113135
rect 335863 113101 335872 113135
rect 335820 113092 335872 113101
rect 244464 113024 244516 113076
rect 261484 111843 261536 111852
rect 261484 111809 261493 111843
rect 261493 111809 261527 111843
rect 261527 111809 261536 111843
rect 261484 111800 261536 111809
rect 331772 111843 331824 111852
rect 331772 111809 331781 111843
rect 331781 111809 331815 111843
rect 331815 111809 331824 111843
rect 331772 111800 331824 111809
rect 232044 111732 232096 111784
rect 232136 111732 232188 111784
rect 334532 111775 334584 111784
rect 334532 111741 334541 111775
rect 334541 111741 334575 111775
rect 334575 111741 334584 111775
rect 334532 111732 334584 111741
rect 317328 109735 317380 109744
rect 317328 109701 317337 109735
rect 317337 109701 317371 109735
rect 317371 109701 317380 109735
rect 317328 109692 317380 109701
rect 344100 109012 344152 109064
rect 344284 109012 344336 109064
rect 3332 108944 3384 108996
rect 31024 108944 31076 108996
rect 340052 108944 340104 108996
rect 253204 108332 253256 108384
rect 317144 107627 317196 107636
rect 317144 107593 317153 107627
rect 317153 107593 317187 107627
rect 317187 107593 317196 107627
rect 317144 107584 317196 107593
rect 232320 107015 232372 107024
rect 232320 106981 232329 107015
rect 232329 106981 232363 107015
rect 232363 106981 232372 107015
rect 232320 106972 232372 106981
rect 244924 106972 244976 107024
rect 245108 106972 245160 107024
rect 297548 106904 297600 106956
rect 100668 106335 100720 106344
rect 100668 106301 100677 106335
rect 100677 106301 100711 106335
rect 100711 106301 100720 106335
rect 100668 106292 100720 106301
rect 231216 106335 231268 106344
rect 231216 106301 231225 106335
rect 231225 106301 231259 106335
rect 231259 106301 231268 106335
rect 231216 106292 231268 106301
rect 258908 106335 258960 106344
rect 258908 106301 258917 106335
rect 258917 106301 258951 106335
rect 258951 106301 258960 106335
rect 258908 106292 258960 106301
rect 260380 106335 260432 106344
rect 260380 106301 260389 106335
rect 260389 106301 260423 106335
rect 260423 106301 260432 106335
rect 260380 106292 260432 106301
rect 317236 106131 317288 106140
rect 317236 106097 317245 106131
rect 317245 106097 317279 106131
rect 317279 106097 317288 106131
rect 317236 106088 317288 106097
rect 321100 106063 321152 106072
rect 321100 106029 321109 106063
rect 321109 106029 321143 106063
rect 321143 106029 321152 106063
rect 321100 106020 321152 106029
rect 246488 104864 246540 104916
rect 246580 104864 246632 104916
rect 254676 104907 254728 104916
rect 254676 104873 254685 104907
rect 254685 104873 254719 104907
rect 254719 104873 254728 104907
rect 254676 104864 254728 104873
rect 263048 104907 263100 104916
rect 263048 104873 263057 104907
rect 263057 104873 263091 104907
rect 263091 104873 263100 104907
rect 263048 104864 263100 104873
rect 316960 104907 317012 104916
rect 316960 104873 316969 104907
rect 316969 104873 317003 104907
rect 317003 104873 317012 104907
rect 316960 104864 317012 104873
rect 322296 104864 322348 104916
rect 322388 104864 322440 104916
rect 107476 104839 107528 104848
rect 107476 104805 107485 104839
rect 107485 104805 107519 104839
rect 107519 104805 107528 104839
rect 107476 104796 107528 104805
rect 244372 103615 244424 103624
rect 244372 103581 244381 103615
rect 244381 103581 244415 103615
rect 244415 103581 244424 103615
rect 244372 103572 244424 103581
rect 261484 103572 261536 103624
rect 261392 103504 261444 103556
rect 294788 103547 294840 103556
rect 294788 103513 294797 103547
rect 294797 103513 294831 103547
rect 294831 103513 294840 103547
rect 294788 103504 294840 103513
rect 295984 103504 296036 103556
rect 296076 103504 296128 103556
rect 321192 103572 321244 103624
rect 329012 103572 329064 103624
rect 330484 103572 330536 103624
rect 335820 103615 335872 103624
rect 335820 103581 335829 103615
rect 335829 103581 335863 103615
rect 335863 103581 335872 103615
rect 335820 103572 335872 103581
rect 326252 103504 326304 103556
rect 328920 103504 328972 103556
rect 330392 103504 330444 103556
rect 244372 103436 244424 103488
rect 244648 103436 244700 103488
rect 253204 103479 253256 103488
rect 253204 103445 253213 103479
rect 253213 103445 253247 103479
rect 253247 103445 253256 103479
rect 253204 103436 253256 103445
rect 258908 103479 258960 103488
rect 258908 103445 258917 103479
rect 258917 103445 258951 103479
rect 258951 103445 258960 103479
rect 258908 103436 258960 103445
rect 263048 103479 263100 103488
rect 263048 103445 263057 103479
rect 263057 103445 263091 103479
rect 263091 103445 263100 103479
rect 263048 103436 263100 103445
rect 264520 103436 264572 103488
rect 265808 103436 265860 103488
rect 293316 103479 293368 103488
rect 293316 103445 293325 103479
rect 293325 103445 293359 103479
rect 293359 103445 293368 103479
rect 293316 103436 293368 103445
rect 319628 103479 319680 103488
rect 319628 103445 319637 103479
rect 319637 103445 319671 103479
rect 319671 103445 319680 103479
rect 319628 103436 319680 103445
rect 321100 103436 321152 103488
rect 321284 103436 321336 103488
rect 322296 103479 322348 103488
rect 322296 103445 322305 103479
rect 322305 103445 322339 103479
rect 322339 103445 322348 103479
rect 322296 103436 322348 103445
rect 331772 103436 331824 103488
rect 331864 103436 331916 103488
rect 333244 103436 333296 103488
rect 333336 103436 333388 103488
rect 335820 103436 335872 103488
rect 321284 103232 321336 103284
rect 334532 102255 334584 102264
rect 334532 102221 334541 102255
rect 334541 102221 334575 102255
rect 334575 102221 334584 102255
rect 334532 102212 334584 102221
rect 298928 102187 298980 102196
rect 298928 102153 298937 102187
rect 298937 102153 298971 102187
rect 298971 102153 298980 102187
rect 298928 102144 298980 102153
rect 300216 102187 300268 102196
rect 300216 102153 300225 102187
rect 300225 102153 300259 102187
rect 300259 102153 300268 102187
rect 300216 102144 300268 102153
rect 301688 102187 301740 102196
rect 301688 102153 301697 102187
rect 301697 102153 301731 102187
rect 301731 102153 301740 102187
rect 301688 102144 301740 102153
rect 232136 102119 232188 102128
rect 232136 102085 232145 102119
rect 232145 102085 232179 102119
rect 232179 102085 232188 102119
rect 232136 102076 232188 102085
rect 328920 102119 328972 102128
rect 328920 102085 328929 102119
rect 328929 102085 328963 102119
rect 328963 102085 328972 102119
rect 328920 102076 328972 102085
rect 334532 102119 334584 102128
rect 334532 102085 334541 102119
rect 334541 102085 334575 102119
rect 334575 102085 334584 102119
rect 334532 102076 334584 102085
rect 297456 100759 297508 100768
rect 297456 100725 297465 100759
rect 297465 100725 297499 100759
rect 297499 100725 297508 100759
rect 297456 100716 297508 100725
rect 261392 99764 261444 99816
rect 232688 99424 232740 99476
rect 246488 99424 246540 99476
rect 231216 99399 231268 99408
rect 231216 99365 231225 99399
rect 231225 99365 231259 99399
rect 231259 99365 231268 99399
rect 231216 99356 231268 99365
rect 244924 99356 244976 99408
rect 232688 99288 232740 99340
rect 245016 99288 245068 99340
rect 231216 96747 231268 96756
rect 231216 96713 231225 96747
rect 231225 96713 231259 96747
rect 231259 96713 231268 96747
rect 231216 96704 231268 96713
rect 297456 96636 297508 96688
rect 345296 96636 345348 96688
rect 345388 96636 345440 96688
rect 100668 96611 100720 96620
rect 100668 96577 100677 96611
rect 100677 96577 100711 96611
rect 100711 96577 100720 96611
rect 100668 96568 100720 96577
rect 297548 96500 297600 96552
rect 107476 95251 107528 95260
rect 107476 95217 107485 95251
rect 107485 95217 107519 95251
rect 107519 95217 107528 95251
rect 107476 95208 107528 95217
rect 254676 95208 254728 95260
rect 254768 95208 254820 95260
rect 294788 95276 294840 95328
rect 246304 95183 246356 95192
rect 246304 95149 246313 95183
rect 246313 95149 246347 95183
rect 246347 95149 246356 95183
rect 246304 95140 246356 95149
rect 253204 95183 253256 95192
rect 253204 95149 253213 95183
rect 253213 95149 253247 95183
rect 253247 95149 253256 95183
rect 253204 95140 253256 95149
rect 257160 95140 257212 95192
rect 265716 95183 265768 95192
rect 265716 95149 265725 95183
rect 265725 95149 265759 95183
rect 265759 95149 265768 95183
rect 265716 95140 265768 95149
rect 294696 95140 294748 95192
rect 340052 95183 340104 95192
rect 340052 95149 340061 95183
rect 340061 95149 340095 95183
rect 340095 95149 340104 95183
rect 340052 95140 340104 95149
rect 232320 93891 232372 93900
rect 232320 93857 232329 93891
rect 232329 93857 232363 93891
rect 232363 93857 232372 93891
rect 232320 93848 232372 93857
rect 258908 93891 258960 93900
rect 258908 93857 258917 93891
rect 258917 93857 258951 93891
rect 258951 93857 258960 93891
rect 258908 93848 258960 93857
rect 263048 93891 263100 93900
rect 263048 93857 263057 93891
rect 263057 93857 263091 93891
rect 263091 93857 263100 93891
rect 263048 93848 263100 93857
rect 264428 93891 264480 93900
rect 264428 93857 264437 93891
rect 264437 93857 264471 93891
rect 264471 93857 264480 93891
rect 264428 93848 264480 93857
rect 293316 93891 293368 93900
rect 293316 93857 293325 93891
rect 293325 93857 293359 93891
rect 293359 93857 293368 93891
rect 293316 93848 293368 93857
rect 295984 93848 296036 93900
rect 296076 93848 296128 93900
rect 319628 93891 319680 93900
rect 319628 93857 319637 93891
rect 319637 93857 319671 93891
rect 319671 93857 319680 93891
rect 319628 93848 319680 93857
rect 321100 93891 321152 93900
rect 321100 93857 321109 93891
rect 321109 93857 321143 93891
rect 321143 93857 321152 93891
rect 321100 93848 321152 93857
rect 322388 93848 322440 93900
rect 330392 93848 330444 93900
rect 330484 93848 330536 93900
rect 335912 93891 335964 93900
rect 335912 93857 335921 93891
rect 335921 93857 335955 93891
rect 335955 93857 335964 93891
rect 335912 93848 335964 93857
rect 298928 93780 298980 93832
rect 300216 93780 300268 93832
rect 301688 93780 301740 93832
rect 299020 93712 299072 93764
rect 300308 93712 300360 93764
rect 301780 93712 301832 93764
rect 232136 92531 232188 92540
rect 232136 92497 232145 92531
rect 232145 92497 232179 92531
rect 232179 92497 232188 92531
rect 232136 92488 232188 92497
rect 329196 92488 329248 92540
rect 334624 92488 334676 92540
rect 263048 89768 263100 89820
rect 232320 89743 232372 89752
rect 232320 89709 232329 89743
rect 232329 89709 232363 89743
rect 232363 89709 232372 89743
rect 232320 89700 232372 89709
rect 344100 89700 344152 89752
rect 344284 89700 344336 89752
rect 263048 89632 263100 89684
rect 296628 89063 296680 89072
rect 296628 89029 296637 89063
rect 296637 89029 296671 89063
rect 296671 89029 296680 89063
rect 296628 89020 296680 89029
rect 379428 87116 379480 87168
rect 386328 87116 386380 87168
rect 100668 87023 100720 87032
rect 100668 86989 100677 87023
rect 100677 86989 100711 87023
rect 100711 86989 100720 87023
rect 100668 86980 100720 86989
rect 246028 86980 246080 87032
rect 249708 86912 249760 86964
rect 252100 86912 252152 86964
rect 246120 86844 246172 86896
rect 296628 86887 296680 86896
rect 296628 86853 296637 86887
rect 296637 86853 296671 86887
rect 296671 86853 296680 86887
rect 296628 86844 296680 86853
rect 253204 85620 253256 85672
rect 244464 85552 244516 85604
rect 244648 85552 244700 85604
rect 246304 85552 246356 85604
rect 246396 85552 246448 85604
rect 257068 85595 257120 85604
rect 257068 85561 257077 85595
rect 257077 85561 257111 85595
rect 257111 85561 257120 85595
rect 257068 85552 257120 85561
rect 260288 85552 260340 85604
rect 260380 85552 260432 85604
rect 264428 85552 264480 85604
rect 264520 85552 264572 85604
rect 265716 85552 265768 85604
rect 265808 85552 265860 85604
rect 294696 85552 294748 85604
rect 294788 85552 294840 85604
rect 322296 85552 322348 85604
rect 322388 85552 322440 85604
rect 331772 85552 331824 85604
rect 331864 85552 331916 85604
rect 333244 85552 333296 85604
rect 333336 85552 333388 85604
rect 340144 85552 340196 85604
rect 107476 85527 107528 85536
rect 107476 85493 107485 85527
rect 107485 85493 107519 85527
rect 107519 85493 107528 85527
rect 107476 85484 107528 85493
rect 261668 85484 261720 85536
rect 232228 85348 232280 85400
rect 232228 85212 232280 85264
rect 321100 84260 321152 84312
rect 253020 84235 253072 84244
rect 253020 84201 253029 84235
rect 253029 84201 253063 84235
rect 253063 84201 253072 84235
rect 253020 84192 253072 84201
rect 258724 84192 258776 84244
rect 258908 84192 258960 84244
rect 244464 84167 244516 84176
rect 244464 84133 244473 84167
rect 244473 84133 244507 84167
rect 244507 84133 244516 84167
rect 244464 84124 244516 84133
rect 245016 84124 245068 84176
rect 245108 84124 245160 84176
rect 261668 84167 261720 84176
rect 261668 84133 261677 84167
rect 261677 84133 261711 84167
rect 261711 84133 261720 84167
rect 261668 84124 261720 84133
rect 264520 84167 264572 84176
rect 264520 84133 264529 84167
rect 264529 84133 264563 84167
rect 264563 84133 264572 84167
rect 264520 84124 264572 84133
rect 265808 84124 265860 84176
rect 266360 84124 266412 84176
rect 293316 84167 293368 84176
rect 293316 84133 293325 84167
rect 293325 84133 293359 84167
rect 293359 84133 293368 84167
rect 293316 84124 293368 84133
rect 294788 84167 294840 84176
rect 294788 84133 294797 84167
rect 294797 84133 294831 84167
rect 294831 84133 294840 84167
rect 294788 84124 294840 84133
rect 319628 84167 319680 84176
rect 319628 84133 319637 84167
rect 319637 84133 319671 84167
rect 319671 84133 319680 84167
rect 319628 84124 319680 84133
rect 326252 84124 326304 84176
rect 326344 84124 326396 84176
rect 253020 84056 253072 84108
rect 253112 84056 253164 84108
rect 263048 83011 263100 83020
rect 263048 82977 263057 83011
rect 263057 82977 263091 83011
rect 263091 82977 263100 83011
rect 263048 82968 263100 82977
rect 320824 82943 320876 82952
rect 320824 82909 320833 82943
rect 320833 82909 320867 82943
rect 320867 82909 320876 82943
rect 320824 82900 320876 82909
rect 320824 82807 320876 82816
rect 320824 82773 320833 82807
rect 320833 82773 320867 82807
rect 320867 82773 320876 82807
rect 320824 82764 320876 82773
rect 329196 82764 329248 82816
rect 232044 81404 232096 81456
rect 232136 81404 232188 81456
rect 231216 80112 231268 80164
rect 243636 80112 243688 80164
rect 231216 79976 231268 80028
rect 243544 79976 243596 80028
rect 246120 77324 246172 77376
rect 100668 77231 100720 77240
rect 100668 77197 100677 77231
rect 100677 77197 100711 77231
rect 100711 77197 100720 77231
rect 100668 77188 100720 77197
rect 243544 77188 243596 77240
rect 243636 77188 243688 77240
rect 244464 77231 244516 77240
rect 244464 77197 244473 77231
rect 244473 77197 244507 77231
rect 244507 77197 244516 77231
rect 244464 77188 244516 77197
rect 314200 77231 314252 77240
rect 314200 77197 314209 77231
rect 314209 77197 314243 77231
rect 314243 77197 314252 77231
rect 314200 77188 314252 77197
rect 317052 77188 317104 77240
rect 318248 77188 318300 77240
rect 314384 77120 314436 77172
rect 317052 77052 317104 77104
rect 314384 76984 314436 77036
rect 107476 75939 107528 75948
rect 107476 75905 107485 75939
rect 107485 75905 107519 75939
rect 107519 75905 107528 75939
rect 107476 75896 107528 75905
rect 232412 75896 232464 75948
rect 258908 75964 258960 76016
rect 260380 75964 260432 76016
rect 333152 75964 333204 76016
rect 331772 75896 331824 75948
rect 254768 75871 254820 75880
rect 254768 75837 254777 75871
rect 254777 75837 254811 75871
rect 254811 75837 254820 75871
rect 254768 75828 254820 75837
rect 258816 75828 258868 75880
rect 260288 75828 260340 75880
rect 333244 75896 333296 75948
rect 341432 75896 341484 75948
rect 341708 75896 341760 75948
rect 331864 75828 331916 75880
rect 333152 75828 333204 75880
rect 333336 75828 333388 75880
rect 322296 74740 322348 74792
rect 261668 74647 261720 74656
rect 261668 74613 261677 74647
rect 261677 74613 261711 74647
rect 261711 74613 261720 74647
rect 261668 74604 261720 74613
rect 322296 74604 322348 74656
rect 246028 74579 246080 74588
rect 246028 74545 246037 74579
rect 246037 74545 246071 74579
rect 246071 74545 246080 74579
rect 246028 74536 246080 74545
rect 253112 74536 253164 74588
rect 257068 74536 257120 74588
rect 257160 74536 257212 74588
rect 264520 74579 264572 74588
rect 264520 74545 264529 74579
rect 264529 74545 264563 74579
rect 264563 74545 264572 74579
rect 293316 74579 293368 74588
rect 264520 74536 264572 74545
rect 293316 74545 293325 74579
rect 293325 74545 293359 74579
rect 293359 74545 293368 74579
rect 293316 74536 293368 74545
rect 294788 74579 294840 74588
rect 294788 74545 294797 74579
rect 294797 74545 294831 74579
rect 294831 74545 294840 74579
rect 294788 74536 294840 74545
rect 295984 74536 296036 74588
rect 296076 74536 296128 74588
rect 319628 74579 319680 74588
rect 319628 74545 319637 74579
rect 319637 74545 319671 74579
rect 319671 74545 319680 74579
rect 319628 74536 319680 74545
rect 265624 74468 265676 74520
rect 265808 74468 265860 74520
rect 322296 74468 322348 74520
rect 253296 74400 253348 74452
rect 322388 74400 322440 74452
rect 321100 73176 321152 73228
rect 253296 73108 253348 73160
rect 232136 73083 232188 73092
rect 232136 73049 232145 73083
rect 232145 73049 232179 73083
rect 232179 73049 232188 73083
rect 232136 73040 232188 73049
rect 329012 71791 329064 71800
rect 329012 71757 329021 71791
rect 329021 71757 329055 71791
rect 329055 71757 329064 71791
rect 329012 71748 329064 71757
rect 254952 69640 255004 69692
rect 100668 67643 100720 67652
rect 100668 67609 100677 67643
rect 100677 67609 100711 67643
rect 100711 67609 100720 67643
rect 100668 67600 100720 67609
rect 231124 67600 231176 67652
rect 231308 67600 231360 67652
rect 232596 67600 232648 67652
rect 232688 67600 232740 67652
rect 263048 67643 263100 67652
rect 263048 67609 263057 67643
rect 263057 67609 263091 67643
rect 263091 67609 263100 67643
rect 263048 67600 263100 67609
rect 314200 67643 314252 67652
rect 314200 67609 314209 67643
rect 314209 67609 314243 67643
rect 314243 67609 314252 67643
rect 314200 67600 314252 67609
rect 316868 67600 316920 67652
rect 316960 67600 317012 67652
rect 318156 67643 318208 67652
rect 318156 67609 318165 67643
rect 318165 67609 318199 67643
rect 318199 67609 318208 67643
rect 318156 67600 318208 67609
rect 345388 67575 345440 67584
rect 345388 67541 345397 67575
rect 345397 67541 345431 67575
rect 345431 67541 345440 67575
rect 345388 67532 345440 67541
rect 260288 66308 260340 66360
rect 260196 66240 260248 66292
rect 330392 66240 330444 66292
rect 330484 66240 330536 66292
rect 331772 66240 331824 66292
rect 331864 66240 331916 66292
rect 333244 66240 333296 66292
rect 333336 66240 333388 66292
rect 334532 66240 334584 66292
rect 334624 66240 334676 66292
rect 335820 66240 335872 66292
rect 335912 66240 335964 66292
rect 107476 66215 107528 66224
rect 107476 66181 107485 66215
rect 107485 66181 107519 66215
rect 107519 66181 107528 66215
rect 107476 66172 107528 66181
rect 231124 66172 231176 66224
rect 231308 66172 231360 66224
rect 232320 66172 232372 66224
rect 232412 66172 232464 66224
rect 314200 66215 314252 66224
rect 314200 66181 314209 66215
rect 314209 66181 314243 66215
rect 314243 66181 314252 66215
rect 314200 66172 314252 66181
rect 258816 64880 258868 64932
rect 258908 64880 258960 64932
rect 260196 64812 260248 64864
rect 260380 64812 260432 64864
rect 264520 64855 264572 64864
rect 264520 64821 264529 64855
rect 264529 64821 264563 64855
rect 264563 64821 264572 64855
rect 264520 64812 264572 64821
rect 265808 64855 265860 64864
rect 265808 64821 265817 64855
rect 265817 64821 265851 64855
rect 265851 64821 265860 64855
rect 265808 64812 265860 64821
rect 293316 64855 293368 64864
rect 293316 64821 293325 64855
rect 293325 64821 293359 64855
rect 293359 64821 293368 64855
rect 293316 64812 293368 64821
rect 294788 64855 294840 64864
rect 294788 64821 294797 64855
rect 294797 64821 294831 64855
rect 294831 64821 294840 64855
rect 294788 64812 294840 64821
rect 319628 64855 319680 64864
rect 319628 64821 319637 64855
rect 319637 64821 319671 64855
rect 319671 64821 319680 64855
rect 319628 64812 319680 64821
rect 322388 64812 322440 64864
rect 253204 63563 253256 63572
rect 253204 63529 253213 63563
rect 253213 63529 253247 63563
rect 253247 63529 253256 63563
rect 253204 63520 253256 63529
rect 254860 63452 254912 63504
rect 321008 63495 321060 63504
rect 321008 63461 321017 63495
rect 321017 63461 321051 63495
rect 321051 63461 321060 63495
rect 321008 63452 321060 63461
rect 326252 63452 326304 63504
rect 326344 63452 326396 63504
rect 331772 63495 331824 63504
rect 331772 63461 331781 63495
rect 331781 63461 331815 63495
rect 331815 63461 331824 63495
rect 331772 63452 331824 63461
rect 334532 61455 334584 61464
rect 334532 61421 334541 61455
rect 334541 61421 334575 61455
rect 334575 61421 334584 61455
rect 334532 61412 334584 61421
rect 258908 60120 258960 60172
rect 258908 59984 258960 60036
rect 296168 59984 296220 60036
rect 244924 57944 244976 57996
rect 245016 57944 245068 57996
rect 345388 57987 345440 57996
rect 345388 57953 345397 57987
rect 345397 57953 345431 57987
rect 345431 57953 345440 57987
rect 345388 57944 345440 57953
rect 100668 57919 100720 57928
rect 100668 57885 100677 57919
rect 100677 57885 100711 57919
rect 100711 57885 100720 57919
rect 100668 57876 100720 57885
rect 246580 57876 246632 57928
rect 107476 56627 107528 56636
rect 107476 56593 107485 56627
rect 107485 56593 107519 56627
rect 107519 56593 107528 56627
rect 107476 56584 107528 56593
rect 314200 56627 314252 56636
rect 314200 56593 314209 56627
rect 314209 56593 314243 56627
rect 314243 56593 314252 56627
rect 314200 56584 314252 56593
rect 240692 56516 240744 56568
rect 244464 56559 244516 56568
rect 244464 56525 244473 56559
rect 244473 56525 244507 56559
rect 244507 56525 244516 56559
rect 244464 56516 244516 56525
rect 261668 55972 261720 56024
rect 265808 55335 265860 55344
rect 265808 55301 265817 55335
rect 265817 55301 265851 55335
rect 265851 55301 265860 55335
rect 265808 55292 265860 55301
rect 322296 55335 322348 55344
rect 322296 55301 322305 55335
rect 322305 55301 322339 55335
rect 322339 55301 322348 55335
rect 322296 55292 322348 55301
rect 231308 55199 231360 55208
rect 231308 55165 231317 55199
rect 231317 55165 231351 55199
rect 231351 55165 231360 55199
rect 231308 55156 231360 55165
rect 265808 55199 265860 55208
rect 265808 55165 265817 55199
rect 265817 55165 265851 55199
rect 265851 55165 265860 55199
rect 265808 55156 265860 55165
rect 299020 55199 299072 55208
rect 299020 55165 299029 55199
rect 299029 55165 299063 55199
rect 299063 55165 299072 55199
rect 299020 55156 299072 55165
rect 300308 55199 300360 55208
rect 300308 55165 300317 55199
rect 300317 55165 300351 55199
rect 300351 55165 300360 55199
rect 300308 55156 300360 55165
rect 301780 55199 301832 55208
rect 301780 55165 301789 55199
rect 301789 55165 301823 55199
rect 301823 55165 301832 55199
rect 301780 55156 301832 55165
rect 322296 55156 322348 55208
rect 322388 55156 322440 55208
rect 254768 53839 254820 53848
rect 254768 53805 254777 53839
rect 254777 53805 254811 53839
rect 254811 53805 254820 53839
rect 254768 53796 254820 53805
rect 331772 53839 331824 53848
rect 331772 53805 331781 53839
rect 331781 53805 331815 53839
rect 331815 53805 331824 53839
rect 331772 53796 331824 53805
rect 326160 52436 326212 52488
rect 326252 52436 326304 52488
rect 329012 52436 329064 52488
rect 329196 52436 329248 52488
rect 333060 51076 333112 51128
rect 340052 51008 340104 51060
rect 340236 51008 340288 51060
rect 333152 50940 333204 50992
rect 253020 50328 253072 50380
rect 253296 50328 253348 50380
rect 345388 48356 345440 48408
rect 100668 48331 100720 48340
rect 100668 48297 100677 48331
rect 100677 48297 100711 48331
rect 100711 48297 100720 48331
rect 100668 48288 100720 48297
rect 244924 48288 244976 48340
rect 245016 48288 245068 48340
rect 246488 48331 246540 48340
rect 246488 48297 246497 48331
rect 246497 48297 246531 48331
rect 246531 48297 246540 48331
rect 246488 48288 246540 48297
rect 344192 48288 344244 48340
rect 344284 48288 344336 48340
rect 345296 48288 345348 48340
rect 257160 47064 257212 47116
rect 240692 46996 240744 47048
rect 232136 46971 232188 46980
rect 232136 46937 232145 46971
rect 232145 46937 232179 46971
rect 232179 46937 232188 46971
rect 232136 46928 232188 46937
rect 244372 46928 244424 46980
rect 257160 46928 257212 46980
rect 261576 46971 261628 46980
rect 261576 46937 261585 46971
rect 261585 46937 261619 46971
rect 261619 46937 261628 46971
rect 261576 46928 261628 46937
rect 264520 46971 264572 46980
rect 264520 46937 264529 46971
rect 264529 46937 264563 46971
rect 264563 46937 264572 46971
rect 264520 46928 264572 46937
rect 293408 46928 293460 46980
rect 294880 46928 294932 46980
rect 296168 46928 296220 46980
rect 319628 46971 319680 46980
rect 319628 46937 319637 46971
rect 319637 46937 319671 46971
rect 319671 46937 319680 46971
rect 319628 46928 319680 46937
rect 334532 46971 334584 46980
rect 334532 46937 334541 46971
rect 334541 46937 334575 46971
rect 334575 46937 334584 46971
rect 334532 46928 334584 46937
rect 341524 46928 341576 46980
rect 341708 46928 341760 46980
rect 107476 46903 107528 46912
rect 107476 46869 107485 46903
rect 107485 46869 107519 46903
rect 107519 46869 107528 46903
rect 107476 46860 107528 46869
rect 240692 46903 240744 46912
rect 240692 46869 240701 46903
rect 240701 46869 240735 46903
rect 240735 46869 240744 46903
rect 240692 46860 240744 46869
rect 314200 46903 314252 46912
rect 314200 46869 314209 46903
rect 314209 46869 314243 46903
rect 314243 46869 314252 46903
rect 314200 46860 314252 46869
rect 231308 45611 231360 45620
rect 231308 45577 231317 45611
rect 231317 45577 231351 45611
rect 231351 45577 231360 45611
rect 231308 45568 231360 45577
rect 265808 45611 265860 45620
rect 265808 45577 265817 45611
rect 265817 45577 265851 45611
rect 265851 45577 265860 45611
rect 265808 45568 265860 45577
rect 299020 45611 299072 45620
rect 299020 45577 299029 45611
rect 299029 45577 299063 45611
rect 299063 45577 299072 45611
rect 299020 45568 299072 45577
rect 300308 45611 300360 45620
rect 300308 45577 300317 45611
rect 300317 45577 300351 45611
rect 300351 45577 300360 45611
rect 300308 45568 300360 45577
rect 301780 45611 301832 45620
rect 301780 45577 301789 45611
rect 301789 45577 301823 45611
rect 301823 45577 301832 45611
rect 301780 45568 301832 45577
rect 321100 45568 321152 45620
rect 253020 45500 253072 45552
rect 254768 45500 254820 45552
rect 257160 45543 257212 45552
rect 257160 45509 257169 45543
rect 257169 45509 257203 45543
rect 257203 45509 257212 45543
rect 257160 45500 257212 45509
rect 264520 45500 264572 45552
rect 319628 45543 319680 45552
rect 319628 45509 319637 45543
rect 319637 45509 319671 45543
rect 319671 45509 319680 45543
rect 319628 45500 319680 45509
rect 322388 45500 322440 45552
rect 254768 45364 254820 45416
rect 326160 44208 326212 44260
rect 326252 44208 326304 44260
rect 329012 44140 329064 44192
rect 329104 44140 329156 44192
rect 326252 44072 326304 44124
rect 331772 44072 331824 44124
rect 331956 44072 332008 44124
rect 261576 42143 261628 42152
rect 261576 42109 261585 42143
rect 261585 42109 261619 42143
rect 261619 42109 261628 42143
rect 261576 42100 261628 42109
rect 244372 41463 244424 41472
rect 244372 41429 244381 41463
rect 244381 41429 244415 41463
rect 244415 41429 244424 41463
rect 244372 41420 244424 41429
rect 344192 41420 344244 41472
rect 344100 41352 344152 41404
rect 232412 40672 232464 40724
rect 232780 40715 232832 40724
rect 232780 40681 232789 40715
rect 232789 40681 232823 40715
rect 232823 40681 232832 40715
rect 232780 40672 232832 40681
rect 252928 40715 252980 40724
rect 252928 40681 252937 40715
rect 252937 40681 252971 40715
rect 252971 40681 252980 40715
rect 252928 40672 252980 40681
rect 321008 40715 321060 40724
rect 321008 40681 321017 40715
rect 321017 40681 321051 40715
rect 321051 40681 321060 40715
rect 321008 40672 321060 40681
rect 322296 40715 322348 40724
rect 322296 40681 322305 40715
rect 322305 40681 322339 40715
rect 322339 40681 322348 40715
rect 322296 40672 322348 40681
rect 335452 40264 335504 40316
rect 344928 40264 344980 40316
rect 345296 38632 345348 38684
rect 345388 38632 345440 38684
rect 100668 38607 100720 38616
rect 100668 38573 100677 38607
rect 100677 38573 100711 38607
rect 100711 38573 100720 38607
rect 100668 38564 100720 38573
rect 244372 38607 244424 38616
rect 244372 38573 244381 38607
rect 244381 38573 244415 38607
rect 244415 38573 244424 38607
rect 244372 38564 244424 38573
rect 240692 37383 240744 37392
rect 240692 37349 240701 37383
rect 240701 37349 240735 37383
rect 240735 37349 240744 37383
rect 240692 37340 240744 37349
rect 265808 37340 265860 37392
rect 107476 37315 107528 37324
rect 107476 37281 107485 37315
rect 107485 37281 107519 37315
rect 107519 37281 107528 37315
rect 107476 37272 107528 37281
rect 258816 37272 258868 37324
rect 258908 37272 258960 37324
rect 314200 37315 314252 37324
rect 314200 37281 314209 37315
rect 314209 37281 314243 37315
rect 314243 37281 314252 37315
rect 314200 37272 314252 37281
rect 240232 37204 240284 37256
rect 240692 37204 240744 37256
rect 261668 35912 261720 35964
rect 264428 35955 264480 35964
rect 264428 35921 264437 35955
rect 264437 35921 264471 35955
rect 264471 35921 264480 35955
rect 264428 35912 264480 35921
rect 265716 35955 265768 35964
rect 265716 35921 265725 35955
rect 265725 35921 265759 35955
rect 265759 35921 265768 35955
rect 265716 35912 265768 35921
rect 319628 35955 319680 35964
rect 319628 35921 319637 35955
rect 319637 35921 319671 35955
rect 319671 35921 319680 35955
rect 319628 35912 319680 35921
rect 252928 35887 252980 35896
rect 252928 35853 252937 35887
rect 252937 35853 252971 35887
rect 252971 35853 252980 35887
rect 252928 35844 252980 35853
rect 299020 35887 299072 35896
rect 299020 35853 299029 35887
rect 299029 35853 299063 35887
rect 299063 35853 299072 35887
rect 299020 35844 299072 35853
rect 300308 35887 300360 35896
rect 300308 35853 300317 35887
rect 300317 35853 300351 35887
rect 300351 35853 300360 35887
rect 300308 35844 300360 35853
rect 301780 35887 301832 35896
rect 301780 35853 301789 35887
rect 301789 35853 301823 35887
rect 301823 35853 301832 35887
rect 301780 35844 301832 35853
rect 245844 33804 245896 33856
rect 246028 33804 246080 33856
rect 262956 31764 263008 31816
rect 319628 31764 319680 31816
rect 319536 31696 319588 31748
rect 321008 31739 321060 31748
rect 321008 31705 321017 31739
rect 321017 31705 321051 31739
rect 321051 31705 321060 31739
rect 321008 31696 321060 31705
rect 263048 31628 263100 31680
rect 379428 29180 379480 29232
rect 386328 29180 386380 29232
rect 240600 29044 240652 29096
rect 100668 29019 100720 29028
rect 100668 28985 100677 29019
rect 100677 28985 100711 29019
rect 100711 28985 100720 29019
rect 100668 28976 100720 28985
rect 264428 28976 264480 29028
rect 264520 28976 264572 29028
rect 265716 28976 265768 29028
rect 265808 28976 265860 29028
rect 267096 28976 267148 29028
rect 267188 28976 267240 29028
rect 268568 28976 268620 29028
rect 268660 28976 268712 29028
rect 333060 28976 333112 29028
rect 240600 28908 240652 28960
rect 244924 28908 244976 28960
rect 245016 28908 245068 28960
rect 340052 28908 340104 28960
rect 333152 28840 333204 28892
rect 339960 28840 340012 28892
rect 232320 27659 232372 27668
rect 232320 27625 232329 27659
rect 232329 27625 232363 27659
rect 232363 27625 232372 27659
rect 232320 27616 232372 27625
rect 232780 27659 232832 27668
rect 232780 27625 232789 27659
rect 232789 27625 232823 27659
rect 232823 27625 232832 27659
rect 232780 27616 232832 27625
rect 257160 27659 257212 27668
rect 257160 27625 257169 27659
rect 257169 27625 257203 27659
rect 257203 27625 257212 27659
rect 257160 27616 257212 27625
rect 326344 27659 326396 27668
rect 326344 27625 326353 27659
rect 326353 27625 326387 27659
rect 326387 27625 326396 27659
rect 326344 27616 326396 27625
rect 107476 27591 107528 27600
rect 107476 27557 107485 27591
rect 107485 27557 107519 27591
rect 107519 27557 107528 27591
rect 107476 27548 107528 27557
rect 244464 27591 244516 27600
rect 244464 27557 244473 27591
rect 244473 27557 244507 27591
rect 244507 27557 244516 27591
rect 244464 27548 244516 27557
rect 314200 27591 314252 27600
rect 314200 27557 314209 27591
rect 314209 27557 314243 27591
rect 314243 27557 314252 27591
rect 314200 27548 314252 27557
rect 253020 26256 253072 26308
rect 299020 26299 299072 26308
rect 299020 26265 299029 26299
rect 299029 26265 299063 26299
rect 299063 26265 299072 26299
rect 299020 26256 299072 26265
rect 300308 26299 300360 26308
rect 300308 26265 300317 26299
rect 300317 26265 300351 26299
rect 300351 26265 300360 26299
rect 300308 26256 300360 26265
rect 301780 26299 301832 26308
rect 301780 26265 301789 26299
rect 301789 26265 301823 26299
rect 301823 26265 301832 26299
rect 301780 26256 301832 26265
rect 329196 24828 329248 24880
rect 329380 24828 329432 24880
rect 297640 23400 297692 23452
rect 297548 23375 297600 23384
rect 297548 23341 297557 23375
rect 297557 23341 297591 23375
rect 297591 23341 297600 23375
rect 297548 23332 297600 23341
rect 2872 22040 2924 22092
rect 349804 22040 349856 22092
rect 326344 19388 326396 19440
rect 237932 19320 237984 19372
rect 238024 19320 238076 19372
rect 242164 19320 242216 19372
rect 242256 19320 242308 19372
rect 243544 19320 243596 19372
rect 243636 19320 243688 19372
rect 245844 19320 245896 19372
rect 246028 19320 246080 19372
rect 326160 19320 326212 19372
rect 344100 19320 344152 19372
rect 344192 19320 344244 19372
rect 345388 19320 345440 19372
rect 345480 19320 345532 19372
rect 100484 19252 100536 19304
rect 100668 19252 100720 19304
rect 110328 19252 110380 19304
rect 346584 19252 346636 19304
rect 103428 19184 103480 19236
rect 345664 19184 345716 19236
rect 99288 19116 99340 19168
rect 343916 19116 343968 19168
rect 96528 19048 96580 19100
rect 342536 19048 342588 19100
rect 92388 18980 92440 19032
rect 342812 18980 342864 19032
rect 89628 18912 89680 18964
rect 341340 18912 341392 18964
rect 85488 18844 85540 18896
rect 341064 18844 341116 18896
rect 82636 18776 82688 18828
rect 339776 18776 339828 18828
rect 78588 18708 78640 18760
rect 339868 18708 339920 18760
rect 74448 18640 74500 18692
rect 338488 18640 338540 18692
rect 5448 18572 5500 18624
rect 324872 18572 324924 18624
rect 294880 18504 294932 18556
rect 443000 18504 443052 18556
rect 301780 18275 301832 18284
rect 301780 18241 301789 18275
rect 301789 18241 301823 18275
rect 301823 18241 301832 18275
rect 301780 18232 301832 18241
rect 301872 18207 301924 18216
rect 301872 18173 301881 18207
rect 301881 18173 301915 18207
rect 301915 18173 301924 18207
rect 301872 18164 301924 18173
rect 304816 18028 304868 18080
rect 322940 18028 322992 18080
rect 332508 18028 332560 18080
rect 240232 17960 240284 18012
rect 240692 17960 240744 18012
rect 244464 18003 244516 18012
rect 244464 17969 244473 18003
rect 244473 17969 244507 18003
rect 244507 17969 244516 18003
rect 244464 17960 244516 17969
rect 246304 17960 246356 18012
rect 246488 17960 246540 18012
rect 304908 18003 304960 18012
rect 304908 17969 304917 18003
rect 304917 17969 304951 18003
rect 304951 17969 304960 18003
rect 304908 17960 304960 17969
rect 314200 18003 314252 18012
rect 314200 17969 314209 18003
rect 314209 17969 314243 18003
rect 314243 17969 314252 18003
rect 314200 17960 314252 17969
rect 329104 18003 329156 18012
rect 329104 17969 329113 18003
rect 329113 17969 329147 18003
rect 329147 17969 329156 18003
rect 329104 17960 329156 17969
rect 293684 17892 293736 17944
rect 431960 17892 432012 17944
rect 253112 17824 253164 17876
rect 253296 17824 253348 17876
rect 293408 17824 293460 17876
rect 433340 17824 433392 17876
rect 293592 17756 293644 17808
rect 434720 17756 434772 17808
rect 293500 17688 293552 17740
rect 436100 17688 436152 17740
rect 294972 17620 295024 17672
rect 438860 17620 438912 17672
rect 295064 17552 295116 17604
rect 440240 17552 440292 17604
rect 303068 17484 303120 17536
rect 483020 17484 483072 17536
rect 304632 17416 304684 17468
rect 485780 17416 485832 17468
rect 304448 17348 304500 17400
rect 485872 17348 485924 17400
rect 302056 17323 302108 17332
rect 302056 17289 302065 17323
rect 302065 17289 302099 17323
rect 302099 17289 302108 17323
rect 302056 17280 302108 17289
rect 304540 17280 304592 17332
rect 488540 17280 488592 17332
rect 301964 17255 302016 17264
rect 301964 17221 301973 17255
rect 301973 17221 302007 17255
rect 302007 17221 302016 17255
rect 301964 17212 302016 17221
rect 302148 17255 302200 17264
rect 302148 17221 302157 17255
rect 302157 17221 302191 17255
rect 302191 17221 302200 17255
rect 302148 17212 302200 17221
rect 304724 17212 304776 17264
rect 489920 17212 489972 17264
rect 278412 17187 278464 17196
rect 278412 17153 278421 17187
rect 278421 17153 278455 17187
rect 278455 17153 278464 17187
rect 278412 17144 278464 17153
rect 278596 17187 278648 17196
rect 278596 17153 278605 17187
rect 278605 17153 278639 17187
rect 278639 17153 278648 17187
rect 278596 17144 278648 17153
rect 285036 17144 285088 17196
rect 390560 17144 390612 17196
rect 278228 17119 278280 17128
rect 278228 17085 278237 17119
rect 278237 17085 278271 17119
rect 278271 17085 278280 17119
rect 278228 17076 278280 17085
rect 278320 17119 278372 17128
rect 278320 17085 278329 17119
rect 278329 17085 278363 17119
rect 278363 17085 278372 17119
rect 278504 17119 278556 17128
rect 278320 17076 278372 17085
rect 278504 17085 278513 17119
rect 278513 17085 278547 17119
rect 278547 17085 278556 17119
rect 278504 17076 278556 17085
rect 278688 17119 278740 17128
rect 278688 17085 278697 17119
rect 278697 17085 278731 17119
rect 278731 17085 278740 17119
rect 278688 17076 278740 17085
rect 283840 17076 283892 17128
rect 387800 17076 387852 17128
rect 274088 17008 274140 17060
rect 339776 17008 339828 17060
rect 274272 16940 274324 16992
rect 339684 16940 339736 16992
rect 274180 16872 274232 16924
rect 336740 16872 336792 16924
rect 505008 16872 505060 16924
rect 511908 16872 511960 16924
rect 272800 16804 272852 16856
rect 335360 16804 335412 16856
rect 272708 16736 272760 16788
rect 332784 16736 332836 16788
rect 268752 16711 268804 16720
rect 268752 16677 268761 16711
rect 268761 16677 268795 16711
rect 268795 16677 268804 16711
rect 268752 16668 268804 16677
rect 268936 16711 268988 16720
rect 268936 16677 268945 16711
rect 268945 16677 268979 16711
rect 268979 16677 268988 16711
rect 268936 16668 268988 16677
rect 272892 16668 272944 16720
rect 331312 16668 331364 16720
rect 394700 16668 394752 16720
rect 404268 16668 404320 16720
rect 268844 16643 268896 16652
rect 268844 16609 268853 16643
rect 268853 16609 268887 16643
rect 268887 16609 268896 16643
rect 268844 16600 268896 16609
rect 269028 16643 269080 16652
rect 269028 16609 269037 16643
rect 269037 16609 269071 16643
rect 269071 16609 269080 16643
rect 269028 16600 269080 16609
rect 272984 16600 273036 16652
rect 330116 16600 330168 16652
rect 330392 16600 330444 16652
rect 330576 16600 330628 16652
rect 331864 16600 331916 16652
rect 331956 16600 332008 16652
rect 437388 16600 437440 16652
rect 442908 16600 442960 16652
rect 67548 16532 67600 16584
rect 337016 16532 337068 16584
rect 64788 16464 64840 16516
rect 337108 16464 337160 16516
rect 60648 16396 60700 16448
rect 335820 16396 335872 16448
rect 56508 16328 56560 16380
rect 335544 16328 335596 16380
rect 53748 16260 53800 16312
rect 334348 16260 334400 16312
rect 49608 16192 49660 16244
rect 334072 16192 334124 16244
rect 345020 16192 345072 16244
rect 346400 16192 346452 16244
rect 45468 16124 45520 16176
rect 332876 16124 332928 16176
rect 41328 16056 41380 16108
rect 331404 16056 331456 16108
rect 38568 15988 38620 16040
rect 331496 15988 331548 16040
rect 34428 15920 34480 15972
rect 330392 15920 330444 15972
rect 30288 15852 30340 15904
rect 330208 15852 330260 15904
rect 95148 15784 95200 15836
rect 342444 15784 342496 15836
rect 99196 15716 99248 15768
rect 343732 15716 343784 15768
rect 102048 15648 102100 15700
rect 344100 15648 344152 15700
rect 106188 15580 106240 15632
rect 345112 15580 345164 15632
rect 108948 15512 109000 15564
rect 345204 15512 345256 15564
rect 113088 15444 113140 15496
rect 346952 15444 347004 15496
rect 117228 15376 117280 15428
rect 348424 15376 348476 15428
rect 119988 15308 120040 15360
rect 348056 15308 348108 15360
rect 124128 15240 124180 15292
rect 349344 15240 349396 15292
rect 301964 15215 302016 15224
rect 301964 15181 301973 15215
rect 301973 15181 302007 15215
rect 302007 15181 302016 15215
rect 301964 15172 302016 15181
rect 302148 15215 302200 15224
rect 302148 15181 302157 15215
rect 302157 15181 302191 15215
rect 302191 15181 302200 15215
rect 302148 15172 302200 15181
rect 304632 15215 304684 15224
rect 304632 15181 304641 15215
rect 304641 15181 304675 15215
rect 304675 15181 304684 15215
rect 304632 15172 304684 15181
rect 304908 15215 304960 15224
rect 304908 15181 304917 15215
rect 304917 15181 304951 15215
rect 304951 15181 304960 15215
rect 304908 15172 304960 15181
rect 307208 15215 307260 15224
rect 307208 15181 307217 15215
rect 307217 15181 307251 15215
rect 307251 15181 307260 15215
rect 307208 15172 307260 15181
rect 329104 15215 329156 15224
rect 329104 15181 329113 15215
rect 329113 15181 329147 15215
rect 329147 15181 329156 15215
rect 329104 15172 329156 15181
rect 302056 15147 302108 15156
rect 302056 15113 302065 15147
rect 302065 15113 302099 15147
rect 302099 15113 302108 15147
rect 302056 15104 302108 15113
rect 303160 15104 303212 15156
rect 477500 15104 477552 15156
rect 303252 15036 303304 15088
rect 481640 15036 481692 15088
rect 91008 14968 91060 15020
rect 342904 14968 342956 15020
rect 88248 14900 88300 14952
rect 340972 14900 341024 14952
rect 84108 14832 84160 14884
rect 341248 14832 341300 14884
rect 81348 14764 81400 14816
rect 339960 14764 340012 14816
rect 77208 14696 77260 14748
rect 339592 14696 339644 14748
rect 73068 14628 73120 14680
rect 338304 14628 338356 14680
rect 70308 14560 70360 14612
rect 338212 14560 338264 14612
rect 66168 14492 66220 14544
rect 336832 14492 336884 14544
rect 63408 14424 63460 14476
rect 337292 14424 337344 14476
rect 474740 14356 474792 14408
rect 470600 14288 470652 14340
rect 300308 14220 300360 14272
rect 467840 14220 467892 14272
rect 300400 14152 300452 14204
rect 463700 14152 463752 14204
rect 299020 14084 299072 14136
rect 459560 14084 459612 14136
rect 456800 14016 456852 14068
rect 452660 13948 452712 14000
rect 296168 13880 296220 13932
rect 449900 13880 449952 13932
rect 296260 13812 296312 13864
rect 445760 13812 445812 13864
rect 281080 13744 281132 13796
rect 374000 13744 374052 13796
rect 283564 13676 283616 13728
rect 378140 13676 378192 13728
rect 282460 13608 282512 13660
rect 382280 13608 382332 13660
rect 283932 13540 283984 13592
rect 385040 13540 385092 13592
rect 284024 13472 284076 13524
rect 389180 13472 389232 13524
rect 285312 13404 285364 13456
rect 391940 13404 391992 13456
rect 285220 13336 285272 13388
rect 396080 13336 396132 13388
rect 286508 13268 286560 13320
rect 400220 13268 400272 13320
rect 287980 13200 288032 13252
rect 402980 13200 403032 13252
rect 268936 13175 268988 13184
rect 268936 13141 268945 13175
rect 268945 13141 268979 13175
rect 268979 13141 268988 13175
rect 268936 13132 268988 13141
rect 287796 13132 287848 13184
rect 407120 13132 407172 13184
rect 268752 13107 268804 13116
rect 268752 13073 268761 13107
rect 268761 13073 268795 13107
rect 268795 13073 268804 13107
rect 268752 13064 268804 13073
rect 269028 13107 269080 13116
rect 269028 13073 269037 13107
rect 269037 13073 269071 13107
rect 269071 13073 269080 13107
rect 269028 13064 269080 13073
rect 278688 13107 278740 13116
rect 278688 13073 278697 13107
rect 278697 13073 278731 13107
rect 278731 13073 278740 13107
rect 278688 13064 278740 13073
rect 289176 13064 289228 13116
rect 409880 13064 409932 13116
rect 280988 12996 281040 13048
rect 371240 12996 371292 13048
rect 279700 12928 279752 12980
rect 367100 12928 367152 12980
rect 279792 12860 279844 12912
rect 364340 12860 364392 12912
rect 360200 12792 360252 12844
rect 356060 12724 356112 12776
rect 276940 12656 276992 12708
rect 353300 12656 353352 12708
rect 276848 12588 276900 12640
rect 349160 12588 349212 12640
rect 268844 12563 268896 12572
rect 268844 12529 268853 12563
rect 268853 12529 268887 12563
rect 268887 12529 268896 12563
rect 268844 12520 268896 12529
rect 275560 12520 275612 12572
rect 346584 12520 346636 12572
rect 244464 12452 244516 12504
rect 244924 12452 244976 12504
rect 274364 12452 274416 12504
rect 342628 12452 342680 12504
rect 244372 12384 244424 12436
rect 244832 12384 244884 12436
rect 275560 12384 275612 12436
rect 275836 12384 275888 12436
rect 307024 12384 307076 12436
rect 307300 12384 307352 12436
rect 308496 12384 308548 12436
rect 308588 12384 308640 12436
rect 309968 12384 310020 12436
rect 310060 12384 310112 12436
rect 520280 12384 520332 12436
rect 311348 12316 311400 12368
rect 312728 12316 312780 12368
rect 524420 12316 524472 12368
rect 312820 12248 312872 12300
rect 528560 12248 528612 12300
rect 314384 12180 314436 12232
rect 531320 12180 531372 12232
rect 314292 12112 314344 12164
rect 535460 12112 535512 12164
rect 278596 12087 278648 12096
rect 278596 12053 278605 12087
rect 278605 12053 278639 12087
rect 278639 12053 278648 12087
rect 278596 12044 278648 12053
rect 315672 12044 315724 12096
rect 538220 12044 538272 12096
rect 315764 11976 315816 12028
rect 542360 11976 542412 12028
rect 317052 11908 317104 11960
rect 546500 11908 546552 11960
rect 316868 11840 316920 11892
rect 549260 11840 549312 11892
rect 318156 11772 318208 11824
rect 553400 11772 553452 11824
rect 318340 11704 318392 11756
rect 556160 11704 556212 11756
rect 311440 11636 311492 11688
rect 517520 11636 517572 11688
rect 309968 11568 310020 11620
rect 513380 11568 513432 11620
rect 308680 11500 308732 11552
rect 510620 11500 510672 11552
rect 308496 11432 308548 11484
rect 506480 11432 506532 11484
rect 502340 11364 502392 11416
rect 307024 11296 307076 11348
rect 499580 11296 499632 11348
rect 306012 11228 306064 11280
rect 495440 11228 495492 11280
rect 271512 11160 271564 11212
rect 328828 11160 328880 11212
rect 271420 11092 271472 11144
rect 324412 11092 324464 11144
rect 314384 11024 314436 11076
rect 314568 11024 314620 11076
rect 322480 11024 322532 11076
rect 322664 11024 322716 11076
rect 345388 11067 345440 11076
rect 345388 11033 345397 11067
rect 345397 11033 345431 11067
rect 345431 11033 345440 11067
rect 345388 11024 345440 11033
rect 292212 10956 292264 11008
rect 426440 10956 426492 11008
rect 293868 10888 293920 10940
rect 430580 10888 430632 10940
rect 293776 10820 293828 10872
rect 433432 10820 433484 10872
rect 295248 10752 295300 10804
rect 437480 10752 437532 10804
rect 295156 10684 295208 10736
rect 441620 10684 441672 10736
rect 296352 10616 296404 10668
rect 444380 10616 444432 10668
rect 296444 10548 296496 10600
rect 448520 10548 448572 10600
rect 297732 10480 297784 10532
rect 451280 10480 451332 10532
rect 297824 10412 297876 10464
rect 455420 10412 455472 10464
rect 299204 10344 299256 10396
rect 459652 10344 459704 10396
rect 299112 10276 299164 10328
rect 462320 10276 462372 10328
rect 292304 10208 292356 10260
rect 423680 10208 423732 10260
rect 290924 10140 290976 10192
rect 419540 10140 419592 10192
rect 289452 10072 289504 10124
rect 416872 10072 416924 10124
rect 289544 10004 289596 10056
rect 412640 10004 412692 10056
rect 288164 9936 288216 9988
rect 408500 9936 408552 9988
rect 288072 9868 288124 9920
rect 405740 9868 405792 9920
rect 288440 9800 288492 9852
rect 401600 9800 401652 9852
rect 286784 9732 286836 9784
rect 398840 9732 398892 9784
rect 107752 9664 107804 9716
rect 232596 9664 232648 9716
rect 232780 9664 232832 9716
rect 267096 9664 267148 9716
rect 267188 9664 267240 9716
rect 268568 9664 268620 9716
rect 268660 9664 268712 9716
rect 285404 9664 285456 9716
rect 394700 9664 394752 9716
rect 91008 9596 91060 9648
rect 100668 9596 100720 9648
rect 108948 9596 109000 9648
rect 359740 9596 359792 9648
rect 363328 9528 363380 9580
rect 167092 9460 167144 9512
rect 237932 9460 237984 9512
rect 279884 9460 279936 9512
rect 366916 9460 366968 9512
rect 169392 9392 169444 9444
rect 239220 9392 239272 9444
rect 281264 9392 281316 9444
rect 370412 9392 370464 9444
rect 165896 9324 165948 9376
rect 237472 9324 237524 9376
rect 281172 9324 281224 9376
rect 374092 9324 374144 9376
rect 164700 9256 164752 9308
rect 237748 9256 237800 9308
rect 282552 9256 282604 9308
rect 377588 9256 377640 9308
rect 163504 9188 163556 9240
rect 237656 9188 237708 9240
rect 282644 9188 282696 9240
rect 381176 9188 381228 9240
rect 162308 9120 162360 9172
rect 236644 9120 236696 9172
rect 268660 9120 268712 9172
rect 314568 9120 314620 9172
rect 161112 9052 161164 9104
rect 236460 9052 236512 9104
rect 270040 9052 270092 9104
rect 318064 9120 318116 9172
rect 318524 9120 318576 9172
rect 317236 9052 317288 9104
rect 545304 9120 545356 9172
rect 129004 8984 129056 9036
rect 230480 8984 230532 9036
rect 271604 8984 271656 9036
rect 324044 9052 324096 9104
rect 552388 9052 552440 9104
rect 577412 8984 577464 9036
rect 126612 8916 126664 8968
rect 229284 8916 229336 8968
rect 269948 8916 270000 8968
rect 321652 8916 321704 8968
rect 322572 8916 322624 8968
rect 324136 8916 324188 8968
rect 581092 8916 581144 8968
rect 277124 8848 277176 8900
rect 356152 8848 356204 8900
rect 277032 8780 277084 8832
rect 352564 8780 352616 8832
rect 275744 8712 275796 8764
rect 349068 8712 349120 8764
rect 275652 8644 275704 8696
rect 345480 8644 345532 8696
rect 274456 8576 274508 8628
rect 341892 8576 341944 8628
rect 274548 8508 274600 8560
rect 338304 8508 338356 8560
rect 273076 8440 273128 8492
rect 334716 8440 334768 8492
rect 273168 8372 273220 8424
rect 331220 8372 331272 8424
rect 271696 8304 271748 8356
rect 327632 8304 327684 8356
rect 328460 8304 328512 8356
rect 328920 8304 328972 8356
rect 345388 8347 345440 8356
rect 345388 8313 345397 8347
rect 345397 8313 345431 8347
rect 345431 8313 345440 8347
rect 345388 8304 345440 8313
rect 196808 8236 196860 8288
rect 244556 8236 244608 8288
rect 252928 8279 252980 8288
rect 252928 8245 252937 8279
rect 252937 8245 252971 8279
rect 252971 8245 252980 8279
rect 252928 8236 252980 8245
rect 302148 8236 302200 8288
rect 472716 8236 472768 8288
rect 193220 8168 193272 8220
rect 243360 8168 243412 8220
rect 302056 8168 302108 8220
rect 476304 8168 476356 8220
rect 189632 8100 189684 8152
rect 243268 8100 243320 8152
rect 303528 8100 303580 8152
rect 479892 8100 479944 8152
rect 186044 8032 186096 8084
rect 241888 8032 241940 8084
rect 304908 8032 304960 8084
rect 484584 8032 484636 8084
rect 182548 7964 182600 8016
rect 241520 7964 241572 8016
rect 304816 7964 304868 8016
rect 488172 7964 488224 8016
rect 178960 7896 179012 7948
rect 240692 7896 240744 7948
rect 264520 7896 264572 7948
rect 293132 7896 293184 7948
rect 306104 7896 306156 7948
rect 491760 7896 491812 7948
rect 175372 7828 175424 7880
rect 239128 7828 239180 7880
rect 265900 7828 265952 7880
rect 296720 7828 296772 7880
rect 306196 7828 306248 7880
rect 495348 7828 495400 7880
rect 171784 7760 171836 7812
rect 239312 7760 239364 7812
rect 265808 7760 265860 7812
rect 300308 7760 300360 7812
rect 307392 7760 307444 7812
rect 307484 7760 307536 7812
rect 498936 7760 498988 7812
rect 168196 7692 168248 7744
rect 237380 7692 237432 7744
rect 267188 7692 267240 7744
rect 303804 7692 303856 7744
rect 502432 7692 502484 7744
rect 157524 7624 157576 7676
rect 236276 7624 236328 7676
rect 267280 7624 267332 7676
rect 307392 7624 307444 7676
rect 308864 7624 308916 7676
rect 506020 7624 506072 7676
rect 153936 7556 153988 7608
rect 234988 7556 235040 7608
rect 268752 7556 268804 7608
rect 310980 7556 311032 7608
rect 311624 7556 311676 7608
rect 520372 7556 520424 7608
rect 200396 7488 200448 7540
rect 244832 7488 244884 7540
rect 300768 7488 300820 7540
rect 469128 7488 469180 7540
rect 203892 7420 203944 7472
rect 246028 7420 246080 7472
rect 300676 7420 300728 7472
rect 465632 7420 465684 7472
rect 207480 7352 207532 7404
rect 246396 7352 246448 7404
rect 299388 7352 299440 7404
rect 462044 7352 462096 7404
rect 211068 7284 211120 7336
rect 247408 7284 247460 7336
rect 299296 7284 299348 7336
rect 458456 7284 458508 7336
rect 214656 7216 214708 7268
rect 247500 7216 247552 7268
rect 297916 7216 297968 7268
rect 454868 7216 454920 7268
rect 218152 7148 218204 7200
rect 248788 7148 248840 7200
rect 298008 7148 298060 7200
rect 451372 7148 451424 7200
rect 221740 7080 221792 7132
rect 248696 7080 248748 7132
rect 296536 7080 296588 7132
rect 447784 7080 447836 7132
rect 225328 7012 225380 7064
rect 250260 7012 250312 7064
rect 296628 7012 296680 7064
rect 444196 7012 444248 7064
rect 228916 6944 228968 6996
rect 250168 6944 250220 6996
rect 270132 6944 270184 6996
rect 320456 6944 320508 6996
rect 322480 6944 322532 6996
rect 328460 6944 328512 6996
rect 331496 6944 331548 6996
rect 332416 6944 332468 6996
rect 339684 6944 339736 6996
rect 340696 6944 340748 6996
rect 329104 6876 329156 6928
rect 329196 6876 329248 6928
rect 332968 6876 333020 6928
rect 333152 6876 333204 6928
rect 195612 6808 195664 6860
rect 243084 6808 243136 6860
rect 281356 6808 281408 6860
rect 376392 6808 376444 6860
rect 192024 6740 192076 6792
rect 243452 6740 243504 6792
rect 260564 6740 260616 6792
rect 271696 6740 271748 6792
rect 282828 6740 282880 6792
rect 379980 6740 380032 6792
rect 188436 6672 188488 6724
rect 242164 6672 242216 6724
rect 258816 6672 258868 6724
rect 269304 6672 269356 6724
rect 282736 6672 282788 6724
rect 383568 6672 383620 6724
rect 184848 6604 184900 6656
rect 241796 6604 241848 6656
rect 260472 6604 260524 6656
rect 272892 6604 272944 6656
rect 284208 6604 284260 6656
rect 387064 6604 387116 6656
rect 181352 6536 181404 6588
rect 240416 6536 240468 6588
rect 261852 6536 261904 6588
rect 276480 6536 276532 6588
rect 285496 6536 285548 6588
rect 390652 6536 390704 6588
rect 177764 6468 177816 6520
rect 240324 6468 240376 6520
rect 260380 6468 260432 6520
rect 275284 6468 275336 6520
rect 285588 6468 285640 6520
rect 394240 6468 394292 6520
rect 174176 6400 174228 6452
rect 238852 6400 238904 6452
rect 261760 6400 261812 6452
rect 278872 6400 278924 6452
rect 286876 6400 286928 6452
rect 397828 6400 397880 6452
rect 170588 6332 170640 6384
rect 238944 6332 238996 6384
rect 261668 6332 261720 6384
rect 286968 6332 287020 6384
rect 401324 6332 401376 6384
rect 159916 6264 159968 6316
rect 236184 6264 236236 6316
rect 261944 6264 261996 6316
rect 282460 6264 282512 6316
rect 288348 6264 288400 6316
rect 404912 6264 404964 6316
rect 156328 6196 156380 6248
rect 236092 6196 236144 6248
rect 262956 6196 263008 6248
rect 285956 6196 286008 6248
rect 288256 6196 288308 6248
rect 408592 6196 408644 6248
rect 152740 6128 152792 6180
rect 235264 6128 235316 6180
rect 263140 6128 263192 6180
rect 289544 6128 289596 6180
rect 289728 6128 289780 6180
rect 412088 6128 412140 6180
rect 199200 6060 199252 6112
rect 244740 6060 244792 6112
rect 281448 6060 281500 6112
rect 372804 6060 372856 6112
rect 202696 5992 202748 6044
rect 245660 5992 245712 6044
rect 279976 5992 280028 6044
rect 369216 5992 369268 6044
rect 206284 5924 206336 5976
rect 245936 5924 245988 5976
rect 280068 5924 280120 5976
rect 365720 5924 365772 5976
rect 209872 5856 209924 5908
rect 247224 5856 247276 5908
rect 278688 5856 278740 5908
rect 362132 5856 362184 5908
rect 213460 5788 213512 5840
rect 247684 5788 247736 5840
rect 278596 5788 278648 5840
rect 358544 5788 358596 5840
rect 217048 5720 217100 5772
rect 248604 5720 248656 5772
rect 277216 5720 277268 5772
rect 354956 5720 355008 5772
rect 220544 5652 220596 5704
rect 248512 5652 248564 5704
rect 277308 5652 277360 5704
rect 351368 5652 351420 5704
rect 224132 5584 224184 5636
rect 250076 5584 250128 5636
rect 275560 5584 275612 5636
rect 347872 5584 347924 5636
rect 227720 5516 227772 5568
rect 249984 5516 250036 5568
rect 252652 5516 252704 5568
rect 275928 5516 275980 5568
rect 344284 5516 344336 5568
rect 124220 5448 124272 5500
rect 191104 5448 191156 5500
rect 194416 5448 194468 5500
rect 243084 5448 243136 5500
rect 243176 5448 243228 5500
rect 254032 5448 254084 5500
rect 255044 5448 255096 5500
rect 255780 5448 255832 5500
rect 256240 5448 256292 5500
rect 257252 5448 257304 5500
rect 257804 5448 257856 5500
rect 258632 5448 258684 5500
rect 264888 5448 264940 5500
rect 291936 5448 291988 5500
rect 311716 5448 311768 5500
rect 522672 5448 522724 5500
rect 113548 5380 113600 5432
rect 182824 5380 182876 5432
rect 187240 5380 187292 5432
rect 241612 5380 241664 5432
rect 241980 5380 242032 5432
rect 257712 5380 257764 5432
rect 259828 5380 259880 5432
rect 264704 5380 264756 5432
rect 294328 5380 294380 5432
rect 313096 5380 313148 5432
rect 526260 5380 526312 5432
rect 125416 5312 125468 5364
rect 195244 5312 195296 5364
rect 198004 5312 198056 5364
rect 244372 5312 244424 5364
rect 244648 5312 244700 5364
rect 254400 5312 254452 5364
rect 257988 5312 258040 5364
rect 261024 5312 261076 5364
rect 264612 5312 264664 5364
rect 267372 5312 267424 5364
rect 295524 5312 295576 5364
rect 313188 5312 313240 5364
rect 529848 5312 529900 5364
rect 158720 5244 158772 5296
rect 235908 5244 235960 5296
rect 236000 5244 236052 5296
rect 251456 5244 251508 5296
rect 257896 5244 257948 5296
rect 262220 5244 262272 5296
rect 266084 5244 266136 5296
rect 297916 5244 297968 5296
rect 314476 5244 314528 5296
rect 533436 5244 533488 5296
rect 155132 5176 155184 5228
rect 235172 5176 235224 5228
rect 238392 5176 238444 5228
rect 252836 5176 252888 5228
rect 266176 5176 266228 5228
rect 299112 5176 299164 5228
rect 314384 5176 314436 5228
rect 536932 5176 536984 5228
rect 151544 5108 151596 5160
rect 234712 5108 234764 5160
rect 237196 5108 237248 5160
rect 252744 5108 252796 5160
rect 266268 5108 266320 5160
rect 301412 5108 301464 5160
rect 315856 5108 315908 5160
rect 540520 5108 540572 5160
rect 148048 5040 148100 5092
rect 233332 5040 233384 5092
rect 234804 5040 234856 5092
rect 251640 5040 251692 5092
rect 267648 5040 267700 5092
rect 144460 4972 144512 5024
rect 233240 4972 233292 5024
rect 233700 4972 233752 5024
rect 251364 4972 251416 5024
rect 260748 4972 260800 5024
rect 270500 4972 270552 5024
rect 302608 5040 302660 5092
rect 315948 5040 316000 5092
rect 544108 5040 544160 5092
rect 305000 4972 305052 5024
rect 317328 4972 317380 5024
rect 547696 4972 547748 5024
rect 140872 4904 140924 4956
rect 232412 4904 232464 4956
rect 232504 4904 232556 4956
rect 251732 4904 251784 4956
rect 259276 4904 259328 4956
rect 268108 4904 268160 4956
rect 306196 4904 306248 4956
rect 318616 4904 318668 4956
rect 551192 4904 551244 4956
rect 133788 4836 133840 4888
rect 231032 4836 231084 4888
rect 231308 4836 231360 4888
rect 251548 4836 251600 4888
rect 262128 4836 262180 4888
rect 267464 4836 267516 4888
rect 308588 4836 308640 4888
rect 318708 4836 318760 4888
rect 554780 4836 554832 4888
rect 127808 4768 127860 4820
rect 229192 4768 229244 4820
rect 230112 4768 230164 4820
rect 251180 4768 251232 4820
rect 262036 4768 262088 4820
rect 265992 4768 266044 4820
rect 106372 4700 106424 4752
rect 120632 4700 120684 4752
rect 186964 4700 187016 4752
rect 201500 4700 201552 4752
rect 244280 4700 244332 4752
rect 245568 4700 245620 4752
rect 254308 4700 254360 4752
rect 260656 4700 260708 4752
rect 268936 4768 268988 4820
rect 312176 4768 312228 4820
rect 320088 4768 320140 4820
rect 558368 4768 558420 4820
rect 290740 4700 290792 4752
rect 311808 4700 311860 4752
rect 519084 4700 519136 4752
rect 172980 4632 173032 4684
rect 239404 4632 239456 4684
rect 239588 4632 239640 4684
rect 252560 4632 252612 4684
rect 263416 4632 263468 4684
rect 287152 4632 287204 4684
rect 310336 4632 310388 4684
rect 515588 4632 515640 4684
rect 180156 4564 180208 4616
rect 238852 4564 238904 4616
rect 173164 4496 173216 4548
rect 208676 4496 208728 4548
rect 212264 4428 212316 4480
rect 238852 4428 238904 4480
rect 240600 4564 240652 4616
rect 240784 4564 240836 4616
rect 246764 4564 246816 4616
rect 254584 4564 254636 4616
rect 263324 4564 263376 4616
rect 288348 4564 288400 4616
rect 310428 4564 310480 4616
rect 512000 4564 512052 4616
rect 247592 4496 247644 4548
rect 247960 4496 248012 4548
rect 254124 4496 254176 4548
rect 259092 4496 259144 4548
rect 263508 4496 263560 4548
rect 284760 4496 284812 4548
rect 309048 4496 309100 4548
rect 508412 4496 508464 4548
rect 246212 4428 246264 4480
rect 250352 4428 250404 4480
rect 255320 4428 255372 4480
rect 263232 4428 263284 4480
rect 283656 4428 283708 4480
rect 308956 4428 309008 4480
rect 504824 4428 504876 4480
rect 215852 4360 215904 4412
rect 247040 4360 247092 4412
rect 251456 4360 251508 4412
rect 255596 4360 255648 4412
rect 259000 4360 259052 4412
rect 263324 4360 263376 4412
rect 180708 4292 180760 4344
rect 219348 4292 219400 4344
rect 222936 4224 222988 4276
rect 249892 4292 249944 4344
rect 252652 4292 252704 4344
rect 255872 4292 255924 4344
rect 259184 4292 259236 4344
rect 226524 4156 226576 4208
rect 248420 4224 248472 4276
rect 249800 4224 249852 4276
rect 253848 4224 253900 4276
rect 255504 4224 255556 4276
rect 281264 4360 281316 4412
rect 307576 4360 307628 4412
rect 501236 4360 501288 4412
rect 265808 4292 265860 4344
rect 277676 4292 277728 4344
rect 307668 4292 307720 4344
rect 497740 4292 497792 4344
rect 267004 4224 267056 4276
rect 274088 4224 274140 4276
rect 292304 4224 292356 4276
rect 306288 4224 306340 4276
rect 494152 4224 494204 4276
rect 249156 4156 249208 4208
rect 254768 4156 254820 4208
rect 259368 4156 259420 4208
rect 264612 4156 264664 4208
rect 264796 4156 264848 4208
rect 271788 4156 271840 4208
rect 326436 4156 326488 4208
rect 330024 4156 330076 4208
rect 36176 4088 36228 4140
rect 37188 4088 37240 4140
rect 37372 4088 37424 4140
rect 38568 4088 38620 4140
rect 42156 4088 42208 4140
rect 42708 4088 42760 4140
rect 44548 4088 44600 4140
rect 45468 4088 45520 4140
rect 55220 4088 55272 4140
rect 56416 4088 56468 4140
rect 334440 4088 334492 4140
rect 46940 4020 46992 4072
rect 332692 4020 332744 4072
rect 45744 3952 45796 4004
rect 332968 3952 333020 4004
rect 39764 3884 39816 3936
rect 331864 3884 331916 3936
rect 38568 3816 38620 3868
rect 180524 3816 180576 3868
rect 263692 3816 263744 3868
rect 331680 3816 331732 3868
rect 32680 3748 32732 3800
rect 329932 3748 329984 3800
rect 31484 3680 31536 3732
rect 27896 3612 27948 3664
rect 12440 3544 12492 3596
rect 13636 3544 13688 3596
rect 26700 3544 26752 3596
rect 27528 3544 27580 3596
rect 33876 3544 33928 3596
rect 34428 3544 34480 3596
rect 93308 3612 93360 3664
rect 93768 3612 93820 3664
rect 94504 3612 94556 3664
rect 95148 3612 95200 3664
rect 95700 3612 95752 3664
rect 96528 3612 96580 3664
rect 98092 3612 98144 3664
rect 99196 3612 99248 3664
rect 101588 3612 101640 3664
rect 102048 3612 102100 3664
rect 102784 3612 102836 3664
rect 103428 3612 103480 3664
rect 105176 3612 105228 3664
rect 106188 3612 106240 3664
rect 112352 3612 112404 3664
rect 113088 3612 113140 3664
rect 114744 3612 114796 3664
rect 115848 3612 115900 3664
rect 115940 3612 115992 3664
rect 117228 3612 117280 3664
rect 119436 3612 119488 3664
rect 119988 3612 120040 3664
rect 121828 3612 121880 3664
rect 122748 3612 122800 3664
rect 123024 3612 123076 3664
rect 124128 3612 124180 3664
rect 180616 3680 180668 3732
rect 180708 3680 180760 3732
rect 273076 3680 273128 3732
rect 273352 3680 273404 3732
rect 292396 3680 292448 3732
rect 292488 3680 292540 3732
rect 224776 3612 224828 3664
rect 224960 3612 225012 3664
rect 263416 3612 263468 3664
rect 292672 3680 292724 3732
rect 311808 3612 311860 3664
rect 313924 3612 313976 3664
rect 316592 3612 316644 3664
rect 282828 3544 282880 3596
rect 316960 3680 317012 3732
rect 324872 3680 324924 3732
rect 328920 3680 328972 3732
rect 337200 3612 337252 3664
rect 433432 3612 433484 3664
rect 434628 3612 434680 3664
rect 477500 3612 477552 3664
rect 478696 3612 478748 3664
rect 485780 3612 485832 3664
rect 486976 3612 487028 3664
rect 572 3476 624 3528
rect 1308 3476 1360 3528
rect 1676 3476 1728 3528
rect 2688 3476 2740 3528
rect 2872 3476 2924 3528
rect 3976 3476 4028 3528
rect 7656 3476 7708 3528
rect 8208 3476 8260 3528
rect 8852 3476 8904 3528
rect 9588 3476 9640 3528
rect 10048 3476 10100 3528
rect 10968 3476 11020 3528
rect 11244 3476 11296 3528
rect 12348 3476 12400 3528
rect 17224 3476 17276 3528
rect 17868 3476 17920 3528
rect 25504 3476 25556 3528
rect 327080 3544 327132 3596
rect 566740 3544 566792 3596
rect 19524 3408 19576 3460
rect 327816 3408 327868 3460
rect 29092 3340 29144 3392
rect 51632 3340 51684 3392
rect 52368 3340 52420 3392
rect 52828 3340 52880 3392
rect 53748 3340 53800 3392
rect 50528 3272 50580 3324
rect 58808 3340 58860 3392
rect 59268 3340 59320 3392
rect 60004 3340 60056 3392
rect 60648 3340 60700 3392
rect 61200 3340 61252 3392
rect 62028 3340 62080 3392
rect 62396 3340 62448 3392
rect 63408 3340 63460 3392
rect 63592 3340 63644 3392
rect 64788 3340 64840 3392
rect 68284 3340 68336 3392
rect 68928 3340 68980 3392
rect 69480 3340 69532 3392
rect 70308 3340 70360 3392
rect 70676 3340 70728 3392
rect 71688 3340 71740 3392
rect 54024 3272 54076 3324
rect 55128 3272 55180 3324
rect 43352 3204 43404 3256
rect 44088 3204 44140 3256
rect 64788 3204 64840 3256
rect 275192 3340 275244 3392
rect 328644 3476 328696 3528
rect 571432 3476 571484 3528
rect 581000 3476 581052 3528
rect 582196 3476 582248 3528
rect 328460 3408 328512 3460
rect 573824 3408 573876 3460
rect 329196 3340 329248 3392
rect 374000 3340 374052 3392
rect 375196 3340 375248 3392
rect 390560 3340 390612 3392
rect 391848 3340 391900 3392
rect 408500 3340 408552 3392
rect 409696 3340 409748 3392
rect 416780 3340 416832 3392
rect 417976 3340 418028 3392
rect 451280 3340 451332 3392
rect 452476 3340 452528 3392
rect 459560 3340 459612 3392
rect 460848 3340 460900 3392
rect 502340 3340 502392 3392
rect 503628 3340 503680 3392
rect 520280 3340 520332 3392
rect 521476 3340 521528 3392
rect 536840 3340 536892 3392
rect 538128 3340 538180 3392
rect 71872 3272 71924 3324
rect 338580 3272 338632 3324
rect 76656 3204 76708 3256
rect 77208 3204 77260 3256
rect 77852 3204 77904 3256
rect 78588 3204 78640 3256
rect 80244 3204 80296 3256
rect 81348 3204 81400 3256
rect 81440 3204 81492 3256
rect 82544 3204 82596 3256
rect 79048 3136 79100 3188
rect 339500 3204 339552 3256
rect 84936 3136 84988 3188
rect 85488 3136 85540 3188
rect 86132 3136 86184 3188
rect 86868 3136 86920 3188
rect 87328 3136 87380 3188
rect 88248 3136 88300 3188
rect 88524 3136 88576 3188
rect 89628 3136 89680 3188
rect 89720 3136 89772 3188
rect 342720 3136 342772 3188
rect 20720 3000 20772 3052
rect 22008 3000 22060 3052
rect 96896 3000 96948 3052
rect 344008 3068 344060 3120
rect 103980 3000 104032 3052
rect 345388 3000 345440 3052
rect 348148 2932 348200 2984
rect 34980 2864 35032 2916
rect 35808 2864 35860 2916
rect 111156 2864 111208 2916
rect 346676 2864 346728 2916
rect 92112 2796 92164 2848
rect 92388 2796 92440 2848
rect 117136 2796 117188 2848
rect 347780 2796 347832 2848
rect 118240 2728 118292 2780
rect 563060 2456 563112 2508
rect 564348 2456 564400 2508
rect 356060 824 356112 876
rect 357348 824 357400 876
rect 5264 552 5316 604
rect 5448 552 5500 604
rect 90916 595 90968 604
rect 90916 561 90925 595
rect 90925 561 90959 595
rect 90959 561 90968 595
rect 90916 552 90968 561
rect 100484 595 100536 604
rect 100484 561 100493 595
rect 100493 561 100527 595
rect 100527 561 100536 595
rect 100484 552 100536 561
rect 107568 552 107620 604
rect 107752 552 107804 604
rect 108764 595 108816 604
rect 108764 561 108773 595
rect 108773 561 108807 595
rect 108807 561 108816 595
rect 108764 552 108816 561
rect 109960 552 110012 604
rect 110328 552 110380 604
rect 280068 595 280120 604
rect 280068 561 280077 595
rect 280077 561 280111 595
rect 280111 561 280120 595
rect 280068 552 280120 561
rect 324412 552 324464 604
rect 325240 552 325292 604
rect 335360 552 335412 604
rect 335912 552 335964 604
rect 336740 552 336792 604
rect 337108 552 337160 604
rect 349160 552 349212 604
rect 350264 552 350316 604
rect 394700 552 394752 604
rect 395436 552 395488 604
rect 401600 552 401652 604
rect 402520 552 402572 604
rect 402980 552 403032 604
rect 403716 552 403768 604
rect 405740 552 405792 604
rect 406108 552 406160 604
rect 409880 552 409932 604
rect 410892 552 410944 604
rect 423680 552 423732 604
rect 423956 552 424008 604
rect 426440 552 426492 604
rect 427544 552 427596 604
rect 427820 552 427872 604
rect 428740 552 428792 604
rect 430580 552 430632 604
rect 431132 552 431184 604
rect 434720 552 434772 604
rect 435824 552 435876 604
rect 436100 552 436152 604
rect 437020 552 437072 604
rect 437480 552 437532 604
rect 438216 552 438268 604
rect 438860 552 438912 604
rect 439412 552 439464 604
rect 452660 552 452712 604
rect 453672 552 453724 604
rect 455420 552 455472 604
rect 456064 552 456116 604
rect 456800 552 456852 604
rect 457260 552 457312 604
rect 462320 552 462372 604
rect 463240 552 463292 604
rect 463700 552 463752 604
rect 464436 552 464488 604
rect 466460 552 466512 604
rect 466828 552 466880 604
rect 469220 552 469272 604
rect 470324 552 470376 604
rect 470600 552 470652 604
rect 471520 552 471572 604
rect 489920 552 489972 604
rect 490564 552 490616 604
rect 495440 552 495492 604
rect 496544 552 496596 604
rect 499580 552 499632 604
rect 500132 552 500184 604
rect 506480 552 506532 604
rect 507216 552 507268 604
rect 510620 552 510672 604
rect 510804 552 510856 604
rect 513380 552 513432 604
rect 514392 552 514444 604
rect 524420 552 524472 604
rect 525064 552 525116 604
rect 538220 552 538272 604
rect 539324 552 539376 604
rect 540980 552 541032 604
rect 541716 552 541768 604
rect 542360 552 542412 604
rect 542912 552 542964 604
rect 549260 552 549312 604
rect 550088 552 550140 604
rect 556160 552 556212 604
rect 557172 552 557224 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700330 8156 703520
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 24320 699718 24348 703520
rect 40512 700398 40540 703520
rect 72988 700534 73016 703520
rect 72976 700528 73028 700534
rect 72976 700470 73028 700476
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 89180 699718 89208 703520
rect 105464 700670 105492 703520
rect 137848 700806 137876 703520
rect 137836 700800 137888 700806
rect 137836 700742 137888 700748
rect 105452 700664 105504 700670
rect 105452 700606 105504 700612
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 89628 699712 89680 699718
rect 89628 699654 89680 699660
rect 3514 682272 3570 682281
rect 3514 682207 3570 682216
rect 3528 681766 3556 682207
rect 3516 681760 3568 681766
rect 3516 681702 3568 681708
rect 3422 667992 3478 668001
rect 3422 667927 3424 667936
rect 3476 667927 3478 667936
rect 3424 667898 3476 667904
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 3422 624880 3478 624889
rect 3422 624815 3478 624824
rect 3436 623830 3464 624815
rect 3424 623824 3476 623830
rect 3424 623766 3476 623772
rect 3422 610464 3478 610473
rect 3422 610399 3478 610408
rect 3436 610026 3464 610399
rect 3424 610020 3476 610026
rect 3424 609962 3476 609968
rect 3238 596048 3294 596057
rect 3238 595983 3294 595992
rect 3252 594862 3280 595983
rect 3240 594856 3292 594862
rect 3240 594798 3292 594804
rect 3422 567352 3478 567361
rect 3422 567287 3478 567296
rect 3436 567254 3464 567287
rect 3424 567248 3476 567254
rect 3424 567190 3476 567196
rect 3146 553072 3202 553081
rect 3146 553007 3202 553016
rect 3160 552090 3188 553007
rect 3148 552084 3200 552090
rect 3148 552026 3200 552032
rect 3422 538656 3478 538665
rect 3422 538591 3478 538600
rect 3436 538286 3464 538591
rect 3424 538280 3476 538286
rect 3424 538222 3476 538228
rect 3422 509960 3478 509969
rect 3422 509895 3478 509904
rect 3436 509386 3464 509895
rect 3424 509380 3476 509386
rect 3424 509322 3476 509328
rect 3422 495544 3478 495553
rect 3422 495479 3424 495488
rect 3476 495479 3478 495488
rect 3424 495450 3476 495456
rect 3146 481128 3202 481137
rect 3146 481063 3202 481072
rect 3160 480282 3188 481063
rect 3148 480276 3200 480282
rect 3148 480218 3200 480224
rect 24780 463078 24808 699654
rect 89640 463146 89668 699654
rect 154132 695570 154160 703520
rect 170324 701010 170352 703520
rect 170312 701004 170364 701010
rect 170312 700946 170364 700952
rect 202800 700194 202828 703520
rect 202788 700188 202840 700194
rect 202788 700130 202840 700136
rect 154120 695564 154172 695570
rect 154120 695506 154172 695512
rect 154212 695564 154264 695570
rect 154212 695506 154264 695512
rect 154224 688634 154252 695506
rect 218992 694210 219020 703520
rect 235184 699990 235212 703520
rect 235172 699984 235224 699990
rect 235172 699926 235224 699932
rect 218980 694204 219032 694210
rect 218980 694146 219032 694152
rect 219164 694204 219216 694210
rect 219164 694146 219216 694152
rect 219176 688702 219204 694146
rect 219164 688696 219216 688702
rect 219164 688638 219216 688644
rect 154212 688628 154264 688634
rect 154212 688570 154264 688576
rect 154396 688628 154448 688634
rect 154396 688570 154448 688576
rect 219072 688628 219124 688634
rect 219072 688570 219124 688576
rect 154408 685846 154436 688570
rect 154396 685840 154448 685846
rect 154396 685782 154448 685788
rect 219084 678994 219112 688570
rect 218992 678966 219112 678994
rect 154304 676252 154356 676258
rect 154304 676194 154356 676200
rect 154316 673538 154344 676194
rect 218992 676190 219020 678966
rect 218980 676184 219032 676190
rect 218980 676126 219032 676132
rect 154304 673532 154356 673538
rect 154304 673474 154356 673480
rect 154488 673532 154540 673538
rect 154488 673474 154540 673480
rect 154500 663762 154528 673474
rect 219072 666596 219124 666602
rect 219072 666538 219124 666544
rect 154316 663734 154528 663762
rect 154316 654158 154344 663734
rect 219084 659682 219112 666538
rect 219084 659666 219204 659682
rect 219084 659660 219216 659666
rect 219084 659654 219164 659660
rect 219164 659602 219216 659608
rect 219348 659660 219400 659666
rect 219348 659602 219400 659608
rect 219360 656878 219388 659602
rect 219348 656872 219400 656878
rect 219348 656814 219400 656820
rect 154304 654152 154356 654158
rect 154304 654094 154356 654100
rect 154488 654152 154540 654158
rect 154488 654094 154540 654100
rect 154500 644450 154528 654094
rect 219256 647284 219308 647290
rect 219256 647226 219308 647232
rect 154316 644422 154528 644450
rect 154316 634846 154344 644422
rect 219268 640422 219296 647226
rect 219256 640416 219308 640422
rect 219256 640358 219308 640364
rect 219072 640280 219124 640286
rect 219072 640222 219124 640228
rect 219084 637566 219112 640222
rect 219072 637560 219124 637566
rect 219072 637502 219124 637508
rect 219164 637560 219216 637566
rect 219164 637502 219216 637508
rect 154304 634840 154356 634846
rect 154304 634782 154356 634788
rect 154488 634840 154540 634846
rect 154488 634782 154540 634788
rect 154500 625138 154528 634782
rect 219176 630578 219204 637502
rect 219176 630550 219388 630578
rect 219360 626550 219388 630550
rect 219348 626544 219400 626550
rect 219348 626486 219400 626492
rect 154316 625110 154528 625138
rect 154316 615534 154344 625110
rect 219348 616888 219400 616894
rect 219348 616830 219400 616836
rect 154304 615528 154356 615534
rect 154304 615470 154356 615476
rect 154488 615528 154540 615534
rect 154488 615470 154540 615476
rect 154500 605826 154528 615470
rect 219360 611454 219388 616830
rect 219348 611448 219400 611454
rect 219348 611390 219400 611396
rect 219072 608728 219124 608734
rect 219072 608670 219124 608676
rect 219084 608598 219112 608670
rect 219072 608592 219124 608598
rect 219072 608534 219124 608540
rect 154316 605798 154528 605826
rect 154316 596222 154344 605798
rect 219256 601588 219308 601594
rect 219256 601530 219308 601536
rect 219268 598942 219296 601530
rect 219256 598936 219308 598942
rect 219256 598878 219308 598884
rect 154304 596216 154356 596222
rect 154488 596216 154540 596222
rect 154304 596158 154356 596164
rect 154408 596164 154488 596170
rect 154408 596158 154540 596164
rect 154408 596142 154528 596158
rect 154408 591954 154436 596142
rect 154316 591926 154436 591954
rect 154316 589286 154344 591926
rect 219164 589348 219216 589354
rect 219164 589290 219216 589296
rect 154304 589280 154356 589286
rect 154304 589222 154356 589228
rect 219176 582418 219204 589290
rect 218980 582412 219032 582418
rect 218980 582354 219032 582360
rect 219164 582412 219216 582418
rect 219164 582354 219216 582360
rect 154304 579760 154356 579766
rect 154224 579708 154304 579714
rect 154224 579702 154356 579708
rect 154224 579686 154344 579702
rect 154224 579630 154252 579686
rect 218992 579630 219020 582354
rect 154212 579624 154264 579630
rect 154212 579566 154264 579572
rect 154396 579624 154448 579630
rect 154396 579566 154448 579572
rect 218980 579624 219032 579630
rect 218980 579566 219032 579572
rect 154408 562970 154436 579566
rect 218888 569968 218940 569974
rect 218888 569910 218940 569916
rect 218900 563106 218928 569910
rect 218888 563100 218940 563106
rect 218888 563042 218940 563048
rect 154212 562964 154264 562970
rect 154212 562906 154264 562912
rect 154396 562964 154448 562970
rect 154396 562906 154448 562912
rect 218980 562964 219032 562970
rect 218980 562906 219032 562912
rect 154224 553330 154252 562906
rect 218992 560266 219020 562906
rect 218900 560238 219020 560266
rect 218900 553450 218928 560238
rect 266268 556232 266320 556238
rect 266268 556174 266320 556180
rect 218888 553444 218940 553450
rect 218888 553386 218940 553392
rect 154224 553302 154344 553330
rect 154316 543810 154344 553302
rect 218888 550656 218940 550662
rect 218888 550598 218940 550604
rect 154316 543782 154528 543810
rect 218900 543794 218928 550598
rect 154500 534018 154528 543782
rect 218888 543788 218940 543794
rect 218888 543730 218940 543736
rect 218980 543652 219032 543658
rect 218980 543594 219032 543600
rect 218992 540977 219020 543594
rect 218978 540968 219034 540977
rect 218978 540903 219034 540912
rect 219162 540968 219218 540977
rect 219162 540903 219218 540912
rect 154408 533990 154528 534018
rect 154408 531282 154436 533990
rect 219176 533882 219204 540903
rect 218992 533854 219204 533882
rect 218992 531321 219020 533854
rect 266176 532772 266228 532778
rect 266176 532714 266228 532720
rect 218978 531312 219034 531321
rect 154396 531276 154448 531282
rect 218978 531247 219034 531256
rect 219162 531312 219218 531321
rect 219162 531247 219218 531256
rect 154396 531218 154448 531224
rect 219176 524346 219204 531247
rect 218980 524340 219032 524346
rect 218980 524282 219032 524288
rect 219164 524340 219216 524346
rect 219164 524282 219216 524288
rect 154488 521688 154540 521694
rect 218992 521665 219020 524282
rect 154488 521630 154540 521636
rect 218794 521656 218850 521665
rect 154500 514706 154528 521630
rect 218794 521591 218850 521600
rect 218978 521656 219034 521665
rect 218978 521591 219034 521600
rect 154408 514678 154528 514706
rect 218808 514690 218836 521591
rect 218796 514684 218848 514690
rect 154408 511970 154436 514678
rect 218796 514626 218848 514632
rect 219072 514684 219124 514690
rect 219072 514626 219124 514632
rect 154396 511964 154448 511970
rect 154396 511906 154448 511912
rect 219084 510610 219112 514626
rect 219072 510604 219124 510610
rect 219072 510546 219124 510552
rect 263508 509312 263560 509318
rect 263508 509254 263560 509260
rect 219072 505096 219124 505102
rect 219072 505038 219124 505044
rect 154488 502376 154540 502382
rect 154488 502318 154540 502324
rect 154500 495394 154528 502318
rect 154316 495366 154528 495394
rect 154316 485858 154344 495366
rect 219084 492726 219112 505038
rect 219072 492720 219124 492726
rect 219072 492662 219124 492668
rect 219164 492720 219216 492726
rect 219164 492662 219216 492668
rect 219176 485858 219204 492662
rect 154304 485852 154356 485858
rect 154304 485794 154356 485800
rect 219164 485852 219216 485858
rect 219164 485794 219216 485800
rect 262128 485852 262180 485858
rect 262128 485794 262180 485800
rect 154396 485716 154448 485722
rect 154396 485658 154448 485664
rect 219256 485716 219308 485722
rect 219256 485658 219308 485664
rect 154408 483002 154436 485658
rect 154396 482996 154448 483002
rect 154396 482938 154448 482944
rect 219268 476134 219296 485658
rect 219072 476128 219124 476134
rect 219072 476070 219124 476076
rect 219256 476128 219308 476134
rect 219256 476070 219308 476076
rect 154396 476060 154448 476066
rect 154396 476002 154448 476008
rect 154408 473362 154436 476002
rect 154408 473334 154528 473362
rect 154500 463729 154528 473334
rect 154302 463720 154358 463729
rect 154302 463655 154358 463664
rect 154486 463720 154542 463729
rect 154486 463655 154542 463664
rect 129752 463406 129872 463434
rect 129752 463350 129780 463406
rect 129740 463344 129792 463350
rect 129740 463286 129792 463292
rect 129844 463282 129872 463406
rect 154316 463350 154344 463655
rect 219084 463418 219112 476070
rect 219072 463412 219124 463418
rect 219072 463354 219124 463360
rect 154304 463344 154356 463350
rect 129832 463276 129884 463282
rect 129832 463218 129884 463224
rect 147692 463270 147812 463298
rect 154304 463286 154356 463292
rect 147692 463214 147720 463270
rect 147680 463208 147732 463214
rect 147680 463150 147732 463156
rect 147784 463146 147812 463270
rect 89628 463140 89680 463146
rect 89628 463082 89680 463088
rect 147772 463140 147824 463146
rect 147772 463082 147824 463088
rect 24768 463072 24820 463078
rect 24768 463014 24820 463020
rect 252466 463040 252522 463049
rect 252466 462975 252522 462984
rect 31024 462936 31076 462942
rect 31024 462878 31076 462884
rect 4620 462868 4672 462874
rect 4620 462810 4672 462816
rect 2964 462800 3016 462806
rect 2964 462742 3016 462748
rect 2780 438048 2832 438054
rect 2778 438016 2780 438025
rect 2832 438016 2834 438025
rect 2778 437951 2834 437960
rect 2976 423745 3004 462742
rect 3240 462732 3292 462738
rect 3240 462674 3292 462680
rect 3148 462664 3200 462670
rect 3148 462606 3200 462612
rect 3056 459400 3108 459406
rect 3056 459342 3108 459348
rect 2962 423736 3018 423745
rect 2962 423671 3018 423680
rect 3068 395049 3096 459342
rect 3054 395040 3110 395049
rect 3054 394975 3110 394984
rect 3160 380633 3188 462606
rect 3146 380624 3202 380633
rect 3146 380559 3202 380568
rect 3252 366217 3280 462674
rect 3424 462392 3476 462398
rect 3424 462334 3476 462340
rect 3330 457736 3386 457745
rect 3330 457671 3386 457680
rect 3238 366208 3294 366217
rect 3238 366143 3294 366152
rect 3344 337521 3372 457671
rect 3330 337512 3386 337521
rect 3330 337447 3386 337456
rect 2780 324216 2832 324222
rect 2780 324158 2832 324164
rect 2792 323105 2820 324158
rect 2778 323096 2834 323105
rect 2778 323031 2834 323040
rect 2780 280152 2832 280158
rect 2778 280120 2780 280129
rect 2832 280120 2834 280129
rect 2778 280055 2834 280064
rect 2780 266144 2832 266150
rect 2780 266086 2832 266092
rect 2792 265713 2820 266086
rect 2778 265704 2834 265713
rect 2778 265639 2834 265648
rect 2780 237312 2832 237318
rect 2780 237254 2832 237260
rect 2792 237017 2820 237254
rect 2778 237008 2834 237017
rect 2778 236943 2834 236952
rect 2780 223100 2832 223106
rect 2780 223042 2832 223048
rect 2792 222601 2820 223042
rect 2778 222592 2834 222601
rect 2778 222527 2834 222536
rect 2780 194336 2832 194342
rect 2780 194278 2832 194284
rect 2792 193905 2820 194278
rect 2778 193896 2834 193905
rect 2778 193831 2834 193840
rect 2780 179716 2832 179722
rect 2780 179658 2832 179664
rect 2792 179489 2820 179658
rect 2778 179480 2834 179489
rect 2778 179415 2834 179424
rect 2780 151360 2832 151366
rect 2780 151302 2832 151308
rect 2792 150793 2820 151302
rect 2778 150784 2834 150793
rect 2778 150719 2834 150728
rect 2780 136400 2832 136406
rect 2778 136368 2780 136377
rect 2832 136368 2834 136377
rect 2778 136303 2834 136312
rect 3332 108996 3384 109002
rect 3332 108938 3384 108944
rect 3344 107681 3372 108938
rect 3330 107672 3386 107681
rect 3330 107607 3386 107616
rect 3330 50960 3386 50969
rect 3330 50895 3386 50904
rect 3344 50153 3372 50895
rect 3330 50144 3386 50153
rect 3330 50079 3386 50088
rect 2872 22092 2924 22098
rect 2872 22034 2924 22040
rect 2884 21457 2912 22034
rect 2870 21448 2926 21457
rect 2870 21383 2926 21392
rect 2686 11792 2742 11801
rect 2686 11727 2742 11736
rect 1306 11656 1362 11665
rect 1306 11591 1362 11600
rect 1320 3534 1348 11591
rect 2700 3534 2728 11727
rect 3436 7177 3464 462334
rect 4068 459332 4120 459338
rect 4068 459274 4120 459280
rect 3976 459196 4028 459202
rect 3976 459138 4028 459144
rect 3884 458992 3936 458998
rect 3884 458934 3936 458940
rect 3792 458924 3844 458930
rect 3792 458866 3844 458872
rect 3700 458720 3752 458726
rect 3700 458662 3752 458668
rect 3608 458448 3660 458454
rect 3608 458390 3660 458396
rect 3516 458380 3568 458386
rect 3516 458322 3568 458328
rect 3528 93265 3556 458322
rect 3620 122097 3648 458390
rect 3712 165073 3740 458662
rect 3804 208185 3832 458866
rect 3896 251297 3924 458934
rect 3988 294409 4016 459138
rect 4080 308825 4108 459274
rect 4632 438054 4660 462810
rect 4712 460216 4764 460222
rect 4712 460158 4764 460164
rect 4620 438048 4672 438054
rect 4620 437990 4672 437996
rect 4724 324222 4752 460158
rect 5448 460148 5500 460154
rect 5448 460090 5500 460096
rect 5264 460080 5316 460086
rect 5264 460022 5316 460028
rect 5080 459944 5132 459950
rect 5080 459886 5132 459892
rect 4896 459808 4948 459814
rect 4896 459750 4948 459756
rect 4804 458652 4856 458658
rect 4804 458594 4856 458600
rect 4712 324216 4764 324222
rect 4712 324158 4764 324164
rect 4066 308816 4122 308825
rect 4066 308751 4122 308760
rect 3974 294400 4030 294409
rect 3974 294335 4030 294344
rect 3882 251288 3938 251297
rect 3882 251223 3938 251232
rect 3790 208176 3846 208185
rect 3790 208111 3846 208120
rect 3698 165064 3754 165073
rect 3698 164999 3754 165008
rect 4816 136406 4844 458594
rect 4908 151366 4936 459750
rect 4988 458788 5040 458794
rect 4988 458730 5040 458736
rect 5000 179722 5028 458730
rect 5092 194342 5120 459886
rect 5172 459060 5224 459066
rect 5172 459002 5224 459008
rect 5184 223106 5212 459002
rect 5276 237318 5304 460022
rect 5356 459128 5408 459134
rect 5356 459070 5408 459076
rect 5368 266150 5396 459070
rect 5460 280158 5488 460090
rect 22006 337648 22062 337657
rect 22006 337583 22062 337592
rect 12346 337512 12402 337521
rect 12346 337447 12402 337456
rect 10966 337376 11022 337385
rect 10966 337311 11022 337320
rect 5448 280152 5500 280158
rect 5448 280094 5500 280100
rect 5356 266144 5408 266150
rect 5356 266086 5408 266092
rect 5264 237312 5316 237318
rect 5264 237254 5316 237260
rect 5172 223100 5224 223106
rect 5172 223042 5224 223048
rect 5080 194336 5132 194342
rect 5080 194278 5132 194284
rect 4988 179716 5040 179722
rect 4988 179658 5040 179664
rect 4896 151360 4948 151366
rect 4896 151302 4948 151308
rect 4804 136400 4856 136406
rect 4804 136342 4856 136348
rect 3606 122088 3662 122097
rect 3606 122023 3662 122032
rect 3514 93256 3570 93265
rect 3514 93191 3570 93200
rect 3514 80064 3570 80073
rect 3514 79999 3570 80008
rect 3528 78985 3556 79999
rect 3514 78976 3570 78985
rect 3514 78911 3570 78920
rect 5448 18624 5500 18630
rect 5448 18566 5500 18572
rect 4066 15872 4122 15881
rect 4066 15807 4122 15816
rect 3974 13016 4030 13025
rect 3974 12951 4030 12960
rect 3422 7168 3478 7177
rect 3422 7103 3478 7112
rect 3988 3534 4016 12951
rect 572 3528 624 3534
rect 572 3470 624 3476
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 1676 3528 1728 3534
rect 1676 3470 1728 3476
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 584 480 612 3470
rect 1688 480 1716 3470
rect 2884 480 2912 3470
rect 4080 480 4108 15807
rect 5460 610 5488 18566
rect 9586 16008 9642 16017
rect 9586 15943 9642 15952
rect 8206 14512 8262 14521
rect 8206 14447 8262 14456
rect 8220 3534 8248 14447
rect 9600 3534 9628 15943
rect 10980 3534 11008 337311
rect 12360 3534 12388 337447
rect 21914 16416 21970 16425
rect 21914 16351 21970 16360
rect 17866 16280 17922 16289
rect 17866 16215 17922 16224
rect 13726 16144 13782 16153
rect 13726 16079 13782 16088
rect 13634 14648 13690 14657
rect 13634 14583 13690 14592
rect 13648 3602 13676 14583
rect 12440 3596 12492 3602
rect 12440 3538 12492 3544
rect 13636 3596 13688 3602
rect 13636 3538 13688 3544
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 12348 3528 12400 3534
rect 12348 3470 12400 3476
rect 6458 3360 6514 3369
rect 6458 3295 6514 3304
rect 5264 604 5316 610
rect 5264 546 5316 552
rect 5448 604 5500 610
rect 5448 546 5500 552
rect 5276 480 5304 546
rect 6472 480 6500 3295
rect 7668 480 7696 3470
rect 8864 480 8892 3470
rect 10060 480 10088 3470
rect 11256 480 11284 3470
rect 12452 480 12480 3538
rect 13740 3482 13768 16079
rect 16026 3632 16082 3641
rect 16026 3567 16082 3576
rect 13648 3454 13768 3482
rect 14830 3496 14886 3505
rect 13648 480 13676 3454
rect 14830 3431 14886 3440
rect 14844 480 14872 3431
rect 16040 480 16068 3567
rect 17880 3534 17908 16215
rect 18326 3768 18382 3777
rect 18326 3703 18382 3712
rect 17224 3528 17276 3534
rect 17224 3470 17276 3476
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 17236 480 17264 3470
rect 18340 480 18368 3703
rect 19524 3460 19576 3466
rect 19524 3402 19576 3408
rect 19536 480 19564 3402
rect 20720 3052 20772 3058
rect 20720 2994 20772 3000
rect 20732 480 20760 2994
rect 21928 480 21956 16351
rect 22020 3058 22048 337583
rect 31036 109002 31064 462878
rect 238760 462528 238812 462534
rect 238760 462470 238812 462476
rect 236644 462460 236696 462466
rect 236644 462402 236696 462408
rect 236656 459884 236684 462402
rect 238772 459884 238800 462470
rect 251638 460048 251694 460057
rect 250720 460012 250772 460018
rect 251638 459983 251694 459992
rect 250720 459954 250772 459960
rect 248326 459912 248382 459921
rect 247250 459882 247632 459898
rect 247250 459876 247644 459882
rect 247250 459870 247592 459876
rect 248262 459870 248326 459898
rect 250732 459898 250760 459954
rect 251652 459898 251680 459983
rect 250378 459870 250760 459898
rect 251390 459870 251680 459898
rect 252480 459884 252508 462975
rect 255594 462768 255650 462777
rect 255594 462703 255650 462712
rect 253478 462496 253534 462505
rect 253478 462431 253534 462440
rect 253492 459884 253520 462431
rect 255608 459884 255636 462703
rect 256606 462632 256662 462641
rect 256606 462567 256662 462576
rect 259828 462596 259880 462602
rect 256620 459884 256648 462567
rect 259828 462538 259880 462544
rect 259840 459884 259868 462538
rect 260840 460284 260892 460290
rect 260840 460226 260892 460232
rect 260852 459884 260880 460226
rect 262140 459898 262168 485794
rect 263520 460034 263548 509254
rect 264888 498228 264940 498234
rect 264888 498170 264940 498176
rect 264900 463010 264928 498170
rect 266188 463010 266216 532714
rect 264060 463004 264112 463010
rect 264060 462946 264112 462952
rect 264888 463004 264940 463010
rect 264888 462946 264940 462952
rect 265072 463004 265124 463010
rect 265072 462946 265124 462952
rect 266176 463004 266228 463010
rect 266176 462946 266228 462952
rect 263244 460006 263548 460034
rect 263244 459898 263272 460006
rect 261970 459870 262168 459898
rect 262982 459870 263272 459898
rect 264072 459884 264100 462946
rect 265084 459884 265112 462946
rect 266280 459898 266308 556174
rect 267556 545148 267608 545154
rect 267556 545090 267608 545096
rect 267568 459898 267596 545090
rect 267660 463486 267688 703520
rect 282828 700732 282880 700738
rect 282828 700674 282880 700680
rect 280068 700460 280120 700466
rect 280068 700402 280120 700408
rect 275928 696992 275980 696998
rect 275928 696934 275980 696940
rect 274548 673532 274600 673538
rect 274548 673474 274600 673480
rect 273168 650072 273220 650078
rect 273168 650014 273220 650020
rect 271788 626612 271840 626618
rect 271788 626554 271840 626560
rect 270408 603152 270460 603158
rect 270408 603094 270460 603100
rect 270316 592068 270368 592074
rect 270316 592010 270368 592016
rect 269028 579692 269080 579698
rect 269028 579634 269080 579640
rect 267648 463480 267700 463486
rect 267648 463422 267700 463428
rect 269040 463010 269068 579634
rect 268200 463004 268252 463010
rect 268200 462946 268252 462952
rect 269028 463004 269080 463010
rect 269028 462946 269080 462952
rect 269304 463004 269356 463010
rect 269304 462946 269356 462952
rect 266110 459870 266308 459898
rect 267214 459870 267596 459898
rect 268212 459884 268240 462946
rect 269316 459884 269344 462946
rect 270328 459884 270356 592010
rect 270420 463010 270448 603094
rect 270408 463004 270460 463010
rect 270408 462946 270460 462952
rect 271800 459898 271828 626554
rect 273180 463010 273208 650014
rect 274456 638988 274508 638994
rect 274456 638930 274508 638936
rect 274468 463010 274496 638930
rect 272432 463004 272484 463010
rect 272432 462946 272484 462952
rect 273168 463004 273220 463010
rect 273168 462946 273220 462952
rect 273444 463004 273496 463010
rect 273444 462946 273496 462952
rect 274456 463004 274508 463010
rect 274456 462946 274508 462952
rect 271446 459870 271828 459898
rect 272444 459884 272472 462946
rect 273456 459884 273484 462946
rect 274560 459884 274588 673474
rect 275940 459898 275968 696934
rect 277308 685908 277360 685914
rect 277308 685850 277360 685856
rect 275586 459870 275968 459898
rect 248326 459847 248382 459856
rect 247592 459818 247644 459824
rect 245382 459776 245438 459785
rect 244030 459746 244136 459762
rect 244030 459740 244148 459746
rect 244030 459734 244096 459740
rect 245134 459734 245382 459762
rect 277320 459762 277348 685850
rect 279792 463208 279844 463214
rect 279792 463150 279844 463156
rect 277676 463140 277728 463146
rect 277676 463082 277728 463088
rect 277688 459884 277716 463082
rect 278780 463004 278832 463010
rect 278780 462946 278832 462952
rect 278792 459884 278820 462946
rect 279804 459884 279832 463150
rect 280080 463010 280108 700402
rect 280896 463548 280948 463554
rect 280896 463490 280948 463496
rect 280068 463004 280120 463010
rect 280068 462946 280120 462952
rect 280908 459884 280936 463490
rect 282840 463214 282868 700674
rect 283852 699854 283880 703520
rect 293224 701004 293276 701010
rect 293224 700946 293276 700952
rect 286968 700936 287020 700942
rect 286968 700878 287020 700884
rect 284208 700868 284260 700874
rect 284208 700810 284260 700816
rect 284116 700596 284168 700602
rect 284116 700538 284168 700544
rect 283840 699848 283892 699854
rect 283840 699790 283892 699796
rect 284128 463214 284156 700538
rect 281908 463208 281960 463214
rect 281908 463150 281960 463156
rect 282828 463208 282880 463214
rect 282828 463150 282880 463156
rect 282920 463208 282972 463214
rect 282920 463150 282972 463156
rect 284116 463208 284168 463214
rect 284116 463150 284168 463156
rect 281920 459884 281948 463150
rect 282932 459884 282960 463150
rect 284220 459898 284248 700810
rect 285588 700256 285640 700262
rect 285588 700198 285640 700204
rect 284050 459870 284248 459898
rect 285600 459762 285628 700198
rect 286980 463214 287008 700878
rect 291844 700188 291896 700194
rect 291844 700130 291896 700136
rect 288348 700120 288400 700126
rect 288348 700062 288400 700068
rect 288256 699916 288308 699922
rect 288256 699858 288308 699864
rect 286140 463208 286192 463214
rect 286140 463150 286192 463156
rect 286968 463208 287020 463214
rect 286968 463150 287020 463156
rect 287152 463208 287204 463214
rect 287152 463150 287204 463156
rect 286152 459884 286180 463150
rect 287164 459884 287192 463150
rect 288268 459884 288296 699858
rect 288360 463214 288388 700062
rect 289728 700052 289780 700058
rect 289728 699994 289780 700000
rect 288348 463208 288400 463214
rect 288348 463150 288400 463156
rect 289740 459762 289768 699994
rect 290464 699984 290516 699990
rect 290464 699926 290516 699932
rect 291108 699984 291160 699990
rect 291108 699926 291160 699932
rect 290476 463622 290504 699926
rect 290464 463616 290516 463622
rect 290464 463558 290516 463564
rect 291120 463214 291148 699926
rect 291292 699848 291344 699854
rect 291292 699790 291344 699796
rect 291304 463842 291332 699790
rect 291304 463814 291608 463842
rect 291384 463684 291436 463690
rect 291384 463626 291436 463632
rect 290372 463208 290424 463214
rect 290372 463150 290424 463156
rect 291108 463208 291160 463214
rect 291108 463150 291160 463156
rect 290384 459884 290412 463150
rect 291396 459884 291424 463626
rect 291580 459898 291608 463814
rect 291856 463690 291884 700130
rect 291844 463684 291896 463690
rect 291844 463626 291896 463632
rect 293236 463418 293264 700946
rect 294604 700800 294656 700806
rect 294604 700742 294656 700748
rect 294512 463684 294564 463690
rect 294512 463626 294564 463632
rect 293500 463616 293552 463622
rect 293500 463558 293552 463564
rect 293224 463412 293276 463418
rect 293224 463354 293276 463360
rect 291580 459870 292422 459898
rect 293512 459884 293540 463558
rect 294524 459884 294552 463626
rect 294616 463350 294644 700742
rect 295984 700664 296036 700670
rect 295984 700606 296036 700612
rect 295996 463486 296024 700606
rect 300136 700534 300164 703520
rect 297364 700528 297416 700534
rect 297364 700470 297416 700476
rect 299480 700528 299532 700534
rect 299480 700470 299532 700476
rect 300124 700528 300176 700534
rect 300124 700470 300176 700476
rect 297376 463690 297404 700470
rect 299492 699990 299520 700470
rect 300124 700392 300176 700398
rect 300124 700334 300176 700340
rect 299480 699984 299532 699990
rect 299480 699926 299532 699932
rect 297364 463684 297416 463690
rect 297364 463626 297416 463632
rect 300136 463622 300164 700334
rect 301504 700324 301556 700330
rect 301504 700266 301556 700272
rect 301516 463690 301544 700266
rect 332520 699922 332548 703520
rect 348804 700058 348832 703520
rect 364996 700126 365024 703520
rect 397472 700262 397500 703520
rect 413664 700942 413692 703520
rect 413652 700936 413704 700942
rect 413652 700878 413704 700884
rect 429856 700874 429884 703520
rect 429844 700868 429896 700874
rect 429844 700810 429896 700816
rect 462332 700738 462360 703520
rect 462320 700732 462372 700738
rect 462320 700674 462372 700680
rect 478524 700602 478552 703520
rect 494808 703474 494836 703520
rect 494808 703446 494928 703474
rect 478512 700596 478564 700602
rect 478512 700538 478564 700544
rect 397460 700256 397512 700262
rect 397460 700198 397512 700204
rect 364984 700120 365036 700126
rect 364984 700062 365036 700068
rect 348792 700052 348844 700058
rect 348792 699994 348844 700000
rect 332508 699916 332560 699922
rect 332508 699858 332560 699864
rect 494900 686089 494928 703446
rect 527192 700466 527220 703520
rect 543476 703474 543504 703520
rect 543476 703446 543596 703474
rect 527180 700460 527232 700466
rect 527180 700402 527232 700408
rect 543568 698290 543596 703446
rect 542728 698284 542780 698290
rect 542728 698226 542780 698232
rect 543556 698284 543608 698290
rect 543556 698226 543608 698232
rect 542740 688702 542768 698226
rect 542728 688696 542780 688702
rect 542728 688638 542780 688644
rect 559668 688634 559696 703520
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 542544 688628 542596 688634
rect 542544 688570 542596 688576
rect 559104 688628 559156 688634
rect 559104 688570 559156 688576
rect 559656 688628 559708 688634
rect 559656 688570 559708 688576
rect 494886 686080 494942 686089
rect 494886 686015 494942 686024
rect 494242 685944 494298 685953
rect 542556 685930 542584 688570
rect 559116 685930 559144 688570
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 494242 685879 494298 685888
rect 542464 685902 542584 685930
rect 559024 685902 559144 685930
rect 580184 685914 580212 686287
rect 580172 685908 580224 685914
rect 305092 681760 305144 681766
rect 305092 681702 305144 681708
rect 300860 463684 300912 463690
rect 300860 463626 300912 463632
rect 301504 463684 301556 463690
rect 301504 463626 301556 463632
rect 303988 463684 304040 463690
rect 303988 463626 304040 463632
rect 298744 463616 298796 463622
rect 298744 463558 298796 463564
rect 300124 463616 300176 463622
rect 300124 463558 300176 463564
rect 295616 463480 295668 463486
rect 295616 463422 295668 463428
rect 295984 463480 296036 463486
rect 295984 463422 296036 463428
rect 294604 463344 294656 463350
rect 294604 463286 294656 463292
rect 295628 459884 295656 463422
rect 296628 463412 296680 463418
rect 296628 463354 296680 463360
rect 296640 459884 296668 463354
rect 297732 463344 297784 463350
rect 297732 463286 297784 463292
rect 297744 459884 297772 463286
rect 298756 459884 298784 463558
rect 299756 463480 299808 463486
rect 299756 463422 299808 463428
rect 299768 459884 299796 463422
rect 300872 459884 300900 463626
rect 302976 463616 303028 463622
rect 302976 463558 303028 463564
rect 301872 463276 301924 463282
rect 301872 463218 301924 463224
rect 301884 459884 301912 463218
rect 302988 459884 303016 463558
rect 304000 459884 304028 463626
rect 305000 463072 305052 463078
rect 305000 463014 305052 463020
rect 305012 459898 305040 463014
rect 305104 460306 305132 681702
rect 494256 678994 494284 685879
rect 542464 684486 542492 685902
rect 559024 684486 559052 685902
rect 580172 685850 580224 685856
rect 542452 684480 542504 684486
rect 542452 684422 542504 684428
rect 559012 684480 559064 684486
rect 559012 684422 559064 684428
rect 494072 678966 494284 678994
rect 494072 676190 494100 678966
rect 494060 676184 494112 676190
rect 494060 676126 494112 676132
rect 580170 674656 580226 674665
rect 580170 674591 580226 674600
rect 580184 673538 580212 674591
rect 580172 673532 580224 673538
rect 580172 673474 580224 673480
rect 305644 667956 305696 667962
rect 305644 667898 305696 667904
rect 305656 463078 305684 667898
rect 494152 666596 494204 666602
rect 494152 666538 494204 666544
rect 542820 666596 542872 666602
rect 542820 666538 542872 666544
rect 559380 666596 559432 666602
rect 559380 666538 559432 666544
rect 494164 659682 494192 666538
rect 542832 659682 542860 666538
rect 559392 659682 559420 666538
rect 494164 659654 494284 659682
rect 494256 654158 494284 659654
rect 542648 659654 542860 659682
rect 559208 659654 559420 659682
rect 494060 654152 494112 654158
rect 494060 654094 494112 654100
rect 494244 654152 494296 654158
rect 494244 654094 494296 654100
rect 306380 652792 306432 652798
rect 306380 652734 306432 652740
rect 305644 463072 305696 463078
rect 305644 463014 305696 463020
rect 305104 460278 305684 460306
rect 305012 459870 305118 459898
rect 276690 459734 277348 459762
rect 285062 459734 285628 459762
rect 289294 459734 289768 459762
rect 305656 459762 305684 460278
rect 306392 460034 306420 652734
rect 494072 644450 494100 654094
rect 542648 647290 542676 659654
rect 559208 647290 559236 659654
rect 580170 651128 580226 651137
rect 580170 651063 580226 651072
rect 580184 650078 580212 651063
rect 580172 650072 580224 650078
rect 580172 650014 580224 650020
rect 542544 647284 542596 647290
rect 542544 647226 542596 647232
rect 542636 647284 542688 647290
rect 542636 647226 542688 647232
rect 559104 647284 559156 647290
rect 559104 647226 559156 647232
rect 559196 647284 559248 647290
rect 559196 647226 559248 647232
rect 494072 644422 494284 644450
rect 494256 634846 494284 644422
rect 542556 640422 542584 647226
rect 559116 640422 559144 647226
rect 542544 640416 542596 640422
rect 542544 640358 542596 640364
rect 542636 640416 542688 640422
rect 542636 640358 542688 640364
rect 559104 640416 559156 640422
rect 559104 640358 559156 640364
rect 559196 640416 559248 640422
rect 559196 640358 559248 640364
rect 494060 634840 494112 634846
rect 494060 634782 494112 634788
rect 494244 634840 494296 634846
rect 494244 634782 494296 634788
rect 494072 625138 494100 634782
rect 542648 630698 542676 640358
rect 559208 630698 559236 640358
rect 580170 639432 580226 639441
rect 580170 639367 580226 639376
rect 580184 638994 580212 639367
rect 580172 638988 580224 638994
rect 580172 638930 580224 638936
rect 542452 630692 542504 630698
rect 542452 630634 542504 630640
rect 542636 630692 542688 630698
rect 542636 630634 542688 630640
rect 559012 630692 559064 630698
rect 559012 630634 559064 630640
rect 559196 630692 559248 630698
rect 559196 630634 559248 630640
rect 542464 630578 542492 630634
rect 559024 630578 559052 630634
rect 542464 630550 542584 630578
rect 559024 630550 559144 630578
rect 494072 625110 494284 625138
rect 309140 623824 309192 623830
rect 309140 623766 309192 623772
rect 308404 610020 308456 610026
rect 308404 609962 308456 609968
rect 308416 463690 308444 609962
rect 308404 463684 308456 463690
rect 308404 463626 308456 463632
rect 308220 463072 308272 463078
rect 308220 463014 308272 463020
rect 306392 460006 306972 460034
rect 306944 459898 306972 460006
rect 306944 459870 307234 459898
rect 308232 459884 308260 463014
rect 309152 459898 309180 623766
rect 494256 615534 494284 625110
rect 542556 621058 542584 630550
rect 559116 621058 559144 630550
rect 580170 627736 580226 627745
rect 580170 627671 580226 627680
rect 580184 626618 580212 627671
rect 580172 626612 580224 626618
rect 580172 626554 580224 626560
rect 542556 621030 542676 621058
rect 559116 621030 559236 621058
rect 494060 615528 494112 615534
rect 494060 615470 494112 615476
rect 494244 615528 494296 615534
rect 494244 615470 494296 615476
rect 494072 605826 494100 615470
rect 542648 611386 542676 621030
rect 559208 611386 559236 621030
rect 542452 611380 542504 611386
rect 542452 611322 542504 611328
rect 542636 611380 542688 611386
rect 542636 611322 542688 611328
rect 559012 611380 559064 611386
rect 559012 611322 559064 611328
rect 559196 611380 559248 611386
rect 559196 611322 559248 611328
rect 542464 611266 542492 611322
rect 559024 611266 559052 611322
rect 542464 611238 542584 611266
rect 559024 611238 559144 611266
rect 542556 608598 542584 611238
rect 559116 608598 559144 611238
rect 542544 608592 542596 608598
rect 542544 608534 542596 608540
rect 559104 608592 559156 608598
rect 559104 608534 559156 608540
rect 494072 605798 494284 605826
rect 494256 596222 494284 605798
rect 580170 604208 580226 604217
rect 580170 604143 580226 604152
rect 580184 603158 580212 604143
rect 580172 603152 580224 603158
rect 580172 603094 580224 603100
rect 542728 601724 542780 601730
rect 542728 601666 542780 601672
rect 559288 601724 559340 601730
rect 559288 601666 559340 601672
rect 542740 598942 542768 601666
rect 559300 598942 559328 601666
rect 542728 598936 542780 598942
rect 542728 598878 542780 598884
rect 559288 598936 559340 598942
rect 559288 598878 559340 598884
rect 494060 596216 494112 596222
rect 494244 596216 494296 596222
rect 494112 596164 494192 596170
rect 494060 596158 494192 596164
rect 494244 596158 494296 596164
rect 494072 596142 494192 596158
rect 494164 596034 494192 596142
rect 494164 596006 494284 596034
rect 309232 594856 309284 594862
rect 309232 594798 309284 594804
rect 309244 460306 309272 594798
rect 494256 591954 494284 596006
rect 580170 592512 580226 592521
rect 580170 592447 580226 592456
rect 580184 592074 580212 592447
rect 580172 592068 580224 592074
rect 580172 592010 580224 592016
rect 494164 591926 494284 591954
rect 494164 589286 494192 591926
rect 542820 589348 542872 589354
rect 542820 589290 542872 589296
rect 559380 589348 559432 589354
rect 559380 589290 559432 589296
rect 493876 589280 493928 589286
rect 493876 589222 493928 589228
rect 494152 589280 494204 589286
rect 494152 589222 494204 589228
rect 493888 579737 493916 589222
rect 542832 582486 542860 589290
rect 559392 582486 559420 589290
rect 542820 582480 542872 582486
rect 542820 582422 542872 582428
rect 559380 582480 559432 582486
rect 559380 582422 559432 582428
rect 542728 582344 542780 582350
rect 542728 582286 542780 582292
rect 559288 582344 559340 582350
rect 559288 582286 559340 582292
rect 493874 579728 493930 579737
rect 493874 579663 493930 579672
rect 494058 579728 494114 579737
rect 494058 579663 494114 579672
rect 494072 572642 494100 579663
rect 542740 572642 542768 582286
rect 559300 572642 559328 582286
rect 580170 580816 580226 580825
rect 580170 580751 580226 580760
rect 580184 579698 580212 580751
rect 580172 579692 580224 579698
rect 580172 579634 580224 579640
rect 494072 572614 494192 572642
rect 494164 569906 494192 572614
rect 542556 572614 542768 572642
rect 559116 572614 559328 572642
rect 542556 569922 542584 572614
rect 559116 569922 559144 572614
rect 494152 569900 494204 569906
rect 494152 569842 494204 569848
rect 542464 569894 542584 569922
rect 559024 569894 559144 569922
rect 311900 567248 311952 567254
rect 311900 567190 311952 567196
rect 311164 552084 311216 552090
rect 311164 552026 311216 552032
rect 311176 463622 311204 552026
rect 311348 463684 311400 463690
rect 311348 463626 311400 463632
rect 311164 463616 311216 463622
rect 311164 463558 311216 463564
rect 309244 460278 309916 460306
rect 309152 459870 309258 459898
rect 309888 459762 309916 460278
rect 311360 459884 311388 463626
rect 311912 460034 311940 567190
rect 542464 563174 542492 569894
rect 559024 563174 559052 569894
rect 542452 563168 542504 563174
rect 542452 563110 542504 563116
rect 559012 563168 559064 563174
rect 559012 563110 559064 563116
rect 494336 563100 494388 563106
rect 494336 563042 494388 563048
rect 494348 560289 494376 563042
rect 542452 563032 542504 563038
rect 542452 562974 542504 562980
rect 559012 563032 559064 563038
rect 559012 562974 559064 562980
rect 494150 560280 494206 560289
rect 494150 560215 494206 560224
rect 494334 560280 494390 560289
rect 542464 560250 542492 562974
rect 559024 560250 559052 562974
rect 494334 560215 494390 560224
rect 542452 560244 542504 560250
rect 494164 550662 494192 560215
rect 542452 560186 542504 560192
rect 559012 560244 559064 560250
rect 559012 560186 559064 560192
rect 580170 557288 580226 557297
rect 580170 557223 580226 557232
rect 580184 556238 580212 557223
rect 580172 556232 580224 556238
rect 580172 556174 580224 556180
rect 494152 550656 494204 550662
rect 494152 550598 494204 550604
rect 494428 550656 494480 550662
rect 494428 550598 494480 550604
rect 542636 550656 542688 550662
rect 542636 550598 542688 550604
rect 559196 550656 559248 550662
rect 559196 550598 559248 550604
rect 494440 543862 494468 550598
rect 494428 543856 494480 543862
rect 494428 543798 494480 543804
rect 494336 543720 494388 543726
rect 494336 543662 494388 543668
rect 494348 540977 494376 543662
rect 542648 543658 542676 550598
rect 559208 543658 559236 550598
rect 580170 545592 580226 545601
rect 580170 545527 580226 545536
rect 580184 545154 580212 545527
rect 580172 545148 580224 545154
rect 580172 545090 580224 545096
rect 542452 543652 542504 543658
rect 542452 543594 542504 543600
rect 542636 543652 542688 543658
rect 542636 543594 542688 543600
rect 559012 543652 559064 543658
rect 559012 543594 559064 543600
rect 559196 543652 559248 543658
rect 559196 543594 559248 543600
rect 494150 540968 494206 540977
rect 494150 540903 494206 540912
rect 494334 540968 494390 540977
rect 494334 540903 494390 540912
rect 313372 538280 313424 538286
rect 313372 538222 313424 538228
rect 311912 460006 312124 460034
rect 312096 459898 312124 460006
rect 313384 459898 313412 538222
rect 494164 531350 494192 540903
rect 542464 534070 542492 543594
rect 559024 534070 559052 543594
rect 542452 534064 542504 534070
rect 542452 534006 542504 534012
rect 542636 534064 542688 534070
rect 542636 534006 542688 534012
rect 559012 534064 559064 534070
rect 559012 534006 559064 534012
rect 559196 534064 559248 534070
rect 559196 534006 559248 534012
rect 494152 531344 494204 531350
rect 494152 531286 494204 531292
rect 494428 531344 494480 531350
rect 494428 531286 494480 531292
rect 494440 524550 494468 531286
rect 494428 524544 494480 524550
rect 494428 524486 494480 524492
rect 542648 524482 542676 534006
rect 559208 524482 559236 534006
rect 580170 533896 580226 533905
rect 580170 533831 580226 533840
rect 580184 532778 580212 533831
rect 580172 532772 580224 532778
rect 580172 532714 580224 532720
rect 542636 524476 542688 524482
rect 542636 524418 542688 524424
rect 559196 524476 559248 524482
rect 559196 524418 559248 524424
rect 494336 524408 494388 524414
rect 494336 524350 494388 524356
rect 542728 524408 542780 524414
rect 542728 524350 542780 524356
rect 559288 524408 559340 524414
rect 559288 524350 559340 524356
rect 494348 521665 494376 524350
rect 542740 521665 542768 524350
rect 559300 521665 559328 524350
rect 494150 521656 494206 521665
rect 494150 521591 494206 521600
rect 494334 521656 494390 521665
rect 494334 521591 494390 521600
rect 542542 521656 542598 521665
rect 542542 521591 542598 521600
rect 542726 521656 542782 521665
rect 542726 521591 542782 521600
rect 559102 521656 559158 521665
rect 559102 521591 559158 521600
rect 559286 521656 559342 521665
rect 559286 521591 559342 521600
rect 494164 512038 494192 521591
rect 542556 512038 542584 521591
rect 559116 512038 559144 521591
rect 494152 512032 494204 512038
rect 494152 511974 494204 511980
rect 494428 512032 494480 512038
rect 494428 511974 494480 511980
rect 542544 512032 542596 512038
rect 542544 511974 542596 511980
rect 542820 512032 542872 512038
rect 542820 511974 542872 511980
rect 559104 512032 559156 512038
rect 559104 511974 559156 511980
rect 559380 512032 559432 512038
rect 559380 511974 559432 511980
rect 314660 509380 314712 509386
rect 314660 509322 314712 509328
rect 313924 495508 313976 495514
rect 313924 495450 313976 495456
rect 313936 463078 313964 495450
rect 314568 463616 314620 463622
rect 314568 463558 314620 463564
rect 313924 463072 313976 463078
rect 313924 463014 313976 463020
rect 312096 459870 312478 459898
rect 313384 459870 313490 459898
rect 314580 459884 314608 463558
rect 314672 460034 314700 509322
rect 494440 502382 494468 511974
rect 542832 502382 542860 511974
rect 559392 502382 559420 511974
rect 580170 510368 580226 510377
rect 580170 510303 580226 510312
rect 580184 509318 580212 510303
rect 580172 509312 580224 509318
rect 580172 509254 580224 509260
rect 494244 502376 494296 502382
rect 493966 502344 494022 502353
rect 493966 502279 494022 502288
rect 494242 502344 494244 502353
rect 494428 502376 494480 502382
rect 494296 502344 494298 502353
rect 542636 502376 542688 502382
rect 494428 502318 494480 502324
rect 542358 502344 542414 502353
rect 494242 502279 494298 502288
rect 542358 502279 542414 502288
rect 542634 502344 542636 502353
rect 542820 502376 542872 502382
rect 542688 502344 542690 502353
rect 559196 502376 559248 502382
rect 542820 502318 542872 502324
rect 558918 502344 558974 502353
rect 542634 502279 542690 502288
rect 558918 502279 558974 502288
rect 559194 502344 559196 502353
rect 559380 502376 559432 502382
rect 559248 502344 559250 502353
rect 559380 502318 559432 502324
rect 559194 502279 559250 502288
rect 493980 492697 494008 502279
rect 542372 492697 542400 502279
rect 558932 492697 558960 502279
rect 580170 498672 580226 498681
rect 580170 498607 580226 498616
rect 580184 498234 580212 498607
rect 580172 498228 580224 498234
rect 580172 498170 580224 498176
rect 493966 492688 494022 492697
rect 493966 492623 494022 492632
rect 494150 492688 494206 492697
rect 494150 492623 494206 492632
rect 542358 492688 542414 492697
rect 542358 492623 542414 492632
rect 542542 492688 542598 492697
rect 542542 492623 542544 492632
rect 494164 489954 494192 492623
rect 542596 492623 542598 492632
rect 558918 492688 558974 492697
rect 558918 492623 558974 492632
rect 559102 492688 559158 492697
rect 559102 492623 559104 492632
rect 542544 492594 542596 492600
rect 559156 492623 559158 492632
rect 559104 492594 559156 492600
rect 494164 489926 494284 489954
rect 494256 480282 494284 489926
rect 580170 486840 580226 486849
rect 580170 486775 580226 486784
rect 580184 485858 580212 486775
rect 580172 485852 580224 485858
rect 580172 485794 580224 485800
rect 542544 485784 542596 485790
rect 542544 485726 542596 485732
rect 559104 485784 559156 485790
rect 559104 485726 559156 485732
rect 542556 483018 542584 485726
rect 559116 483018 559144 485726
rect 542556 482990 542676 483018
rect 559116 482990 559236 483018
rect 316040 480276 316092 480282
rect 316040 480218 316092 480224
rect 494060 480276 494112 480282
rect 494060 480218 494112 480224
rect 494244 480276 494296 480282
rect 494244 480218 494296 480224
rect 314672 460006 315252 460034
rect 315224 459898 315252 460006
rect 315224 459870 315606 459898
rect 316052 459762 316080 480218
rect 494072 480162 494100 480218
rect 494072 480134 494192 480162
rect 494164 470642 494192 480134
rect 542648 476134 542676 482990
rect 559208 476134 559236 482990
rect 542452 476128 542504 476134
rect 542636 476128 542688 476134
rect 542504 476076 542636 476082
rect 542452 476070 542688 476076
rect 559012 476128 559064 476134
rect 559196 476128 559248 476134
rect 559064 476076 559196 476082
rect 559012 476070 559248 476076
rect 542464 476054 542676 476070
rect 559024 476054 559236 476070
rect 494164 470614 494284 470642
rect 494256 463214 494284 470614
rect 542648 466546 542676 476054
rect 559208 466546 559236 476054
rect 542636 466540 542688 466546
rect 542636 466482 542688 466488
rect 559196 466540 559248 466546
rect 559196 466482 559248 466488
rect 542544 463752 542596 463758
rect 542544 463694 542596 463700
rect 559104 463752 559156 463758
rect 559104 463694 559156 463700
rect 494244 463208 494296 463214
rect 494244 463150 494296 463156
rect 542556 463146 542584 463694
rect 542544 463140 542596 463146
rect 542544 463082 542596 463088
rect 317696 463072 317748 463078
rect 317696 463014 317748 463020
rect 317708 459884 317736 463014
rect 559116 463010 559144 463694
rect 580078 463448 580134 463457
rect 580078 463383 580134 463392
rect 559104 463004 559156 463010
rect 559104 462946 559156 462952
rect 342904 462936 342956 462942
rect 318706 462904 318762 462913
rect 342904 462878 342956 462884
rect 318706 462839 318762 462848
rect 320824 462868 320876 462874
rect 318720 459884 318748 462839
rect 320824 462810 320876 462816
rect 319812 462800 319864 462806
rect 319812 462742 319864 462748
rect 319824 459884 319852 462742
rect 320836 459884 320864 462810
rect 322940 462732 322992 462738
rect 322940 462674 322992 462680
rect 322952 459884 322980 462674
rect 324044 462664 324096 462670
rect 324044 462606 324096 462612
rect 324056 459884 324084 462606
rect 327172 460216 327224 460222
rect 327172 460158 327224 460164
rect 327184 459884 327212 460158
rect 330300 460148 330352 460154
rect 330300 460090 330352 460096
rect 330312 459884 330340 460090
rect 333060 460080 333112 460086
rect 333060 460022 333112 460028
rect 333072 459898 333100 460022
rect 336372 459944 336424 459950
rect 333072 459870 333454 459898
rect 336424 459892 336674 459898
rect 336372 459886 336674 459892
rect 336384 459870 336674 459886
rect 342916 459884 342944 462878
rect 580092 462602 580120 463383
rect 580080 462596 580132 462602
rect 580080 462538 580132 462544
rect 577504 462528 577556 462534
rect 577504 462470 577556 462476
rect 348240 462392 348292 462398
rect 348240 462334 348292 462340
rect 348252 459884 348280 462334
rect 339500 459808 339552 459814
rect 305656 459734 306130 459762
rect 309888 459734 310362 459762
rect 316052 459734 316618 459762
rect 339552 459756 339802 459762
rect 339500 459750 339802 459756
rect 339512 459734 339802 459750
rect 245382 459711 245438 459720
rect 244096 459682 244148 459688
rect 241152 459672 241204 459678
rect 231674 459640 231730 459649
rect 231426 459598 231674 459626
rect 232686 459640 232742 459649
rect 232438 459598 232686 459626
rect 231674 459575 231730 459584
rect 233790 459640 233846 459649
rect 233542 459598 233790 459626
rect 232686 459575 232742 459584
rect 235658 459610 235948 459626
rect 240902 459620 241152 459626
rect 242254 459640 242310 459649
rect 240902 459614 241204 459620
rect 235658 459604 235960 459610
rect 235658 459598 235908 459604
rect 233790 459575 233846 459584
rect 240902 459598 241192 459614
rect 241914 459598 242254 459626
rect 242254 459575 242310 459584
rect 343730 459640 343786 459649
rect 345294 459640 345350 459649
rect 343786 459598 344034 459626
rect 345046 459598 345294 459626
rect 343730 459575 343786 459584
rect 345294 459575 345350 459584
rect 235908 459546 235960 459552
rect 237774 459474 238064 459490
rect 239798 459474 240088 459490
rect 243018 459474 243400 459490
rect 246146 459474 246528 459490
rect 249274 459474 249656 459490
rect 254610 459474 254992 459490
rect 257738 459474 258028 459490
rect 237774 459468 238076 459474
rect 237774 459462 238024 459468
rect 239798 459468 240100 459474
rect 239798 459462 240048 459468
rect 238024 459410 238076 459416
rect 243018 459468 243412 459474
rect 243018 459462 243360 459468
rect 240048 459410 240100 459416
rect 246146 459468 246540 459474
rect 246146 459462 246488 459468
rect 243360 459410 243412 459416
rect 249274 459468 249668 459474
rect 249274 459462 249616 459468
rect 246488 459410 246540 459416
rect 254610 459468 255004 459474
rect 254610 459462 254952 459468
rect 249616 459410 249668 459416
rect 257738 459468 258040 459474
rect 257738 459462 257988 459468
rect 254952 459410 255004 459416
rect 257988 459410 258040 459416
rect 349896 459468 349948 459474
rect 349896 459410 349948 459416
rect 321652 459400 321704 459406
rect 234342 459368 234398 459377
rect 229112 459326 230414 459354
rect 86868 338088 86920 338094
rect 86868 338030 86920 338036
rect 82728 337952 82780 337958
rect 82728 337894 82780 337900
rect 75828 337884 75880 337890
rect 75828 337826 75880 337832
rect 62028 337816 62080 337822
rect 37186 337784 37242 337793
rect 62028 337758 62080 337764
rect 37186 337719 37242 337728
rect 35808 337408 35860 337414
rect 35808 337350 35860 337356
rect 31024 108996 31076 109002
rect 31024 108938 31076 108944
rect 27526 16552 27582 16561
rect 27526 16487 27582 16496
rect 24306 4040 24362 4049
rect 24306 3975 24362 3984
rect 23110 3904 23166 3913
rect 23110 3839 23166 3848
rect 22008 3052 22060 3058
rect 22008 2994 22060 3000
rect 23124 480 23152 3839
rect 24320 480 24348 3975
rect 27540 3602 27568 16487
rect 34428 15972 34480 15978
rect 34428 15914 34480 15920
rect 30288 15904 30340 15910
rect 30288 15846 30340 15852
rect 27896 3664 27948 3670
rect 27896 3606 27948 3612
rect 26700 3596 26752 3602
rect 26700 3538 26752 3544
rect 27528 3596 27580 3602
rect 27528 3538 27580 3544
rect 25504 3528 25556 3534
rect 25504 3470 25556 3476
rect 25516 480 25544 3470
rect 26712 480 26740 3538
rect 27908 480 27936 3606
rect 29092 3392 29144 3398
rect 29092 3334 29144 3340
rect 29104 480 29132 3334
rect 30300 480 30328 15846
rect 32680 3800 32732 3806
rect 32680 3742 32732 3748
rect 31484 3732 31536 3738
rect 31484 3674 31536 3680
rect 31496 480 31524 3674
rect 32692 480 32720 3742
rect 34440 3602 34468 15914
rect 33876 3596 33928 3602
rect 33876 3538 33928 3544
rect 34428 3596 34480 3602
rect 34428 3538 34480 3544
rect 33888 480 33916 3538
rect 35820 2922 35848 337350
rect 37200 4146 37228 337719
rect 57888 337680 57940 337686
rect 57888 337622 57940 337628
rect 44088 337612 44140 337618
rect 44088 337554 44140 337560
rect 42708 337476 42760 337482
rect 42708 337418 42760 337424
rect 41328 16108 41380 16114
rect 41328 16050 41380 16056
rect 38568 16040 38620 16046
rect 38568 15982 38620 15988
rect 38580 4146 38608 15982
rect 41340 4842 41368 16050
rect 40972 4814 41368 4842
rect 36176 4140 36228 4146
rect 36176 4082 36228 4088
rect 37188 4140 37240 4146
rect 37188 4082 37240 4088
rect 37372 4140 37424 4146
rect 37372 4082 37424 4088
rect 38568 4140 38620 4146
rect 38568 4082 38620 4088
rect 34980 2916 35032 2922
rect 34980 2858 35032 2864
rect 35808 2916 35860 2922
rect 35808 2858 35860 2864
rect 34992 480 35020 2858
rect 36188 480 36216 4082
rect 37384 480 37412 4082
rect 39764 3936 39816 3942
rect 39764 3878 39816 3884
rect 38568 3868 38620 3874
rect 38568 3810 38620 3816
rect 38580 480 38608 3810
rect 39776 480 39804 3878
rect 40972 480 41000 4814
rect 42720 4146 42748 337418
rect 42156 4140 42208 4146
rect 42156 4082 42208 4088
rect 42708 4140 42760 4146
rect 42708 4082 42760 4088
rect 42168 480 42196 4082
rect 44100 3262 44128 337554
rect 55128 337544 55180 337550
rect 55128 337486 55180 337492
rect 53748 16312 53800 16318
rect 53748 16254 53800 16260
rect 49608 16244 49660 16250
rect 49608 16186 49660 16192
rect 45468 16176 45520 16182
rect 45468 16118 45520 16124
rect 45480 4146 45508 16118
rect 48226 14784 48282 14793
rect 48226 14719 48282 14728
rect 44548 4140 44600 4146
rect 44548 4082 44600 4088
rect 45468 4140 45520 4146
rect 45468 4082 45520 4088
rect 43352 3256 43404 3262
rect 43352 3198 43404 3204
rect 44088 3256 44140 3262
rect 44088 3198 44140 3204
rect 43364 480 43392 3198
rect 44560 480 44588 4082
rect 46940 4072 46992 4078
rect 46940 4014 46992 4020
rect 45744 4004 45796 4010
rect 45744 3946 45796 3952
rect 45756 480 45784 3946
rect 46952 480 46980 4014
rect 48240 3482 48268 14719
rect 49620 3482 49648 16186
rect 52366 14920 52422 14929
rect 52366 14855 52422 14864
rect 48148 3454 48268 3482
rect 49344 3454 49648 3482
rect 48148 480 48176 3454
rect 49344 480 49372 3454
rect 52380 3398 52408 14855
rect 53760 3398 53788 16254
rect 51632 3392 51684 3398
rect 51632 3334 51684 3340
rect 52368 3392 52420 3398
rect 52368 3334 52420 3340
rect 52828 3392 52880 3398
rect 52828 3334 52880 3340
rect 53748 3392 53800 3398
rect 53748 3334 53800 3340
rect 50528 3324 50580 3330
rect 50528 3266 50580 3272
rect 50540 480 50568 3266
rect 51644 480 51672 3334
rect 52840 480 52868 3334
rect 55140 3330 55168 337486
rect 56508 16380 56560 16386
rect 56508 16322 56560 16328
rect 56414 15056 56470 15065
rect 56414 14991 56470 15000
rect 56428 4146 56456 14991
rect 55220 4140 55272 4146
rect 55220 4082 55272 4088
rect 56416 4140 56468 4146
rect 56416 4082 56468 4088
rect 54024 3324 54076 3330
rect 54024 3266 54076 3272
rect 55128 3324 55180 3330
rect 55128 3266 55180 3272
rect 54036 480 54064 3266
rect 55232 480 55260 4082
rect 56520 3482 56548 16322
rect 56428 3454 56548 3482
rect 56428 480 56456 3454
rect 57900 626 57928 337622
rect 60648 16448 60700 16454
rect 60648 16390 60700 16396
rect 59266 15192 59322 15201
rect 59266 15127 59322 15136
rect 59280 3398 59308 15127
rect 60660 3398 60688 16390
rect 62040 3398 62068 337758
rect 68928 337748 68980 337754
rect 68928 337690 68980 337696
rect 67548 16584 67600 16590
rect 67548 16526 67600 16532
rect 64788 16516 64840 16522
rect 64788 16458 64840 16464
rect 63408 14476 63460 14482
rect 63408 14418 63460 14424
rect 63420 3398 63448 14418
rect 64800 3398 64828 16458
rect 66168 14544 66220 14550
rect 66168 14486 66220 14492
rect 66180 3482 66208 14486
rect 67560 3482 67588 16526
rect 65996 3454 66208 3482
rect 67192 3454 67588 3482
rect 58808 3392 58860 3398
rect 58808 3334 58860 3340
rect 59268 3392 59320 3398
rect 59268 3334 59320 3340
rect 60004 3392 60056 3398
rect 60004 3334 60056 3340
rect 60648 3392 60700 3398
rect 60648 3334 60700 3340
rect 61200 3392 61252 3398
rect 61200 3334 61252 3340
rect 62028 3392 62080 3398
rect 62028 3334 62080 3340
rect 62396 3392 62448 3398
rect 62396 3334 62448 3340
rect 63408 3392 63460 3398
rect 63408 3334 63460 3340
rect 63592 3392 63644 3398
rect 63592 3334 63644 3340
rect 64788 3392 64840 3398
rect 64788 3334 64840 3340
rect 57624 598 57928 626
rect 57624 480 57652 598
rect 58820 480 58848 3334
rect 60016 480 60044 3334
rect 61212 480 61240 3334
rect 62408 480 62436 3334
rect 63604 480 63632 3334
rect 64788 3256 64840 3262
rect 64788 3198 64840 3204
rect 64800 480 64828 3198
rect 65996 480 66024 3454
rect 67192 480 67220 3454
rect 68940 3398 68968 337690
rect 74448 18692 74500 18698
rect 74448 18634 74500 18640
rect 71686 17232 71742 17241
rect 71686 17167 71742 17176
rect 70308 14612 70360 14618
rect 70308 14554 70360 14560
rect 70320 3398 70348 14554
rect 71700 3398 71728 17167
rect 73068 14680 73120 14686
rect 73068 14622 73120 14628
rect 68284 3392 68336 3398
rect 68284 3334 68336 3340
rect 68928 3392 68980 3398
rect 68928 3334 68980 3340
rect 69480 3392 69532 3398
rect 69480 3334 69532 3340
rect 70308 3392 70360 3398
rect 70308 3334 70360 3340
rect 70676 3392 70728 3398
rect 70676 3334 70728 3340
rect 71688 3392 71740 3398
rect 71688 3334 71740 3340
rect 68296 480 68324 3334
rect 69492 480 69520 3334
rect 70688 480 70716 3334
rect 71872 3324 71924 3330
rect 71872 3266 71924 3272
rect 71884 480 71912 3266
rect 73080 480 73108 14622
rect 74460 3482 74488 18634
rect 75840 3482 75868 337826
rect 82636 18828 82688 18834
rect 82636 18770 82688 18776
rect 78588 18760 78640 18766
rect 78588 18702 78640 18708
rect 77208 14748 77260 14754
rect 77208 14690 77260 14696
rect 74276 3454 74488 3482
rect 75472 3454 75868 3482
rect 74276 480 74304 3454
rect 75472 480 75500 3454
rect 77220 3262 77248 14690
rect 78600 3262 78628 18702
rect 81348 14816 81400 14822
rect 81348 14758 81400 14764
rect 81360 3262 81388 14758
rect 82648 3618 82676 18770
rect 82556 3590 82676 3618
rect 82556 3262 82584 3590
rect 82740 3482 82768 337894
rect 85488 18896 85540 18902
rect 85488 18838 85540 18844
rect 84108 14884 84160 14890
rect 84108 14826 84160 14832
rect 84120 3482 84148 14826
rect 82648 3454 82768 3482
rect 83844 3454 84148 3482
rect 76656 3256 76708 3262
rect 76656 3198 76708 3204
rect 77208 3256 77260 3262
rect 77208 3198 77260 3204
rect 77852 3256 77904 3262
rect 77852 3198 77904 3204
rect 78588 3256 78640 3262
rect 78588 3198 78640 3204
rect 80244 3256 80296 3262
rect 80244 3198 80296 3204
rect 81348 3256 81400 3262
rect 81348 3198 81400 3204
rect 81440 3256 81492 3262
rect 81440 3198 81492 3204
rect 82544 3256 82596 3262
rect 82544 3198 82596 3204
rect 76668 480 76696 3198
rect 77864 480 77892 3198
rect 79048 3188 79100 3194
rect 79048 3130 79100 3136
rect 79060 480 79088 3130
rect 80256 480 80284 3198
rect 81452 480 81480 3198
rect 82648 480 82676 3454
rect 83844 480 83872 3454
rect 85500 3194 85528 18838
rect 86880 3194 86908 338030
rect 93768 338020 93820 338026
rect 93768 337962 93820 337968
rect 92388 19032 92440 19038
rect 92388 18974 92440 18980
rect 89628 18964 89680 18970
rect 89628 18906 89680 18912
rect 88248 14952 88300 14958
rect 88248 14894 88300 14900
rect 88260 3194 88288 14894
rect 89640 3194 89668 18906
rect 91008 15020 91060 15026
rect 91008 14962 91060 14968
rect 91020 9654 91048 14962
rect 91008 9648 91060 9654
rect 91008 9590 91060 9596
rect 84936 3188 84988 3194
rect 84936 3130 84988 3136
rect 85488 3188 85540 3194
rect 85488 3130 85540 3136
rect 86132 3188 86184 3194
rect 86132 3130 86184 3136
rect 86868 3188 86920 3194
rect 86868 3130 86920 3136
rect 87328 3188 87380 3194
rect 87328 3130 87380 3136
rect 88248 3188 88300 3194
rect 88248 3130 88300 3136
rect 88524 3188 88576 3194
rect 88524 3130 88576 3136
rect 89628 3188 89680 3194
rect 89628 3130 89680 3136
rect 89720 3188 89772 3194
rect 89720 3130 89772 3136
rect 84948 480 84976 3130
rect 86144 480 86172 3130
rect 87340 480 87368 3130
rect 88536 480 88564 3130
rect 89732 480 89760 3130
rect 92400 2854 92428 18974
rect 93780 3670 93808 337962
rect 100668 337340 100720 337346
rect 100668 337282 100720 337288
rect 100680 328438 100708 337282
rect 107476 337272 107528 337278
rect 107476 337214 107528 337220
rect 107488 336734 107516 337214
rect 115848 337204 115900 337210
rect 115848 337146 115900 337152
rect 107476 336728 107528 336734
rect 107476 336670 107528 336676
rect 100668 328432 100720 328438
rect 100668 328374 100720 328380
rect 107476 327140 107528 327146
rect 107476 327082 107528 327088
rect 100668 318844 100720 318850
rect 100668 318786 100720 318792
rect 100680 309126 100708 318786
rect 107488 317422 107516 327082
rect 107476 317416 107528 317422
rect 107476 317358 107528 317364
rect 100668 309120 100720 309126
rect 100668 309062 100720 309068
rect 107476 307828 107528 307834
rect 107476 307770 107528 307776
rect 100668 299532 100720 299538
rect 100668 299474 100720 299480
rect 100680 289814 100708 299474
rect 107488 298110 107516 307770
rect 107476 298104 107528 298110
rect 107476 298046 107528 298052
rect 100668 289808 100720 289814
rect 100668 289750 100720 289756
rect 107476 288448 107528 288454
rect 107476 288390 107528 288396
rect 100668 280220 100720 280226
rect 100668 280162 100720 280168
rect 100680 270502 100708 280162
rect 107488 278769 107516 288390
rect 107474 278760 107530 278769
rect 107474 278695 107530 278704
rect 107658 278760 107714 278769
rect 107658 278695 107714 278704
rect 100668 270496 100720 270502
rect 100668 270438 100720 270444
rect 107672 269142 107700 278695
rect 107476 269136 107528 269142
rect 107476 269078 107528 269084
rect 107660 269136 107712 269142
rect 107660 269078 107712 269084
rect 100668 260908 100720 260914
rect 100668 260850 100720 260856
rect 100680 251190 100708 260850
rect 107488 259457 107516 269078
rect 107474 259448 107530 259457
rect 107474 259383 107530 259392
rect 107658 259448 107714 259457
rect 107658 259383 107714 259392
rect 100668 251184 100720 251190
rect 100668 251126 100720 251132
rect 107672 249830 107700 259383
rect 107476 249824 107528 249830
rect 107476 249766 107528 249772
rect 107660 249824 107712 249830
rect 107660 249766 107712 249772
rect 107488 241777 107516 249766
rect 107474 241768 107530 241777
rect 107474 241703 107530 241712
rect 107474 241632 107530 241641
rect 107474 241567 107530 241576
rect 100668 241528 100720 241534
rect 100668 241470 100720 241476
rect 100680 231849 100708 241470
rect 107488 240145 107516 241567
rect 107474 240136 107530 240145
rect 107474 240071 107530 240080
rect 107658 240136 107714 240145
rect 107658 240071 107714 240080
rect 100666 231840 100722 231849
rect 100666 231775 100722 231784
rect 100850 231840 100906 231849
rect 100850 231775 100906 231784
rect 100864 222222 100892 231775
rect 107672 230518 107700 240071
rect 107476 230512 107528 230518
rect 107476 230454 107528 230460
rect 107660 230512 107712 230518
rect 107660 230454 107712 230460
rect 100668 222216 100720 222222
rect 100668 222158 100720 222164
rect 100852 222216 100904 222222
rect 100852 222158 100904 222164
rect 100680 212537 100708 222158
rect 107488 220833 107516 230454
rect 107474 220824 107530 220833
rect 107474 220759 107530 220768
rect 107658 220824 107714 220833
rect 107658 220759 107714 220768
rect 100666 212528 100722 212537
rect 100666 212463 100722 212472
rect 100850 212528 100906 212537
rect 100850 212463 100906 212472
rect 100864 202910 100892 212463
rect 107672 211177 107700 220759
rect 107474 211168 107530 211177
rect 107474 211103 107530 211112
rect 107658 211168 107714 211177
rect 107658 211103 107714 211112
rect 100668 202904 100720 202910
rect 100668 202846 100720 202852
rect 100852 202904 100904 202910
rect 100852 202846 100904 202852
rect 100680 193225 100708 202846
rect 107488 201482 107516 211103
rect 107476 201476 107528 201482
rect 107476 201418 107528 201424
rect 107660 201476 107712 201482
rect 107660 201418 107712 201424
rect 100666 193216 100722 193225
rect 100666 193151 100722 193160
rect 100850 193216 100906 193225
rect 100850 193151 100906 193160
rect 100864 183598 100892 193151
rect 107672 191865 107700 201418
rect 107474 191856 107530 191865
rect 107474 191791 107530 191800
rect 107658 191856 107714 191865
rect 107658 191791 107714 191800
rect 100668 183592 100720 183598
rect 100668 183534 100720 183540
rect 100852 183592 100904 183598
rect 100852 183534 100904 183540
rect 100680 173913 100708 183534
rect 107488 182170 107516 191791
rect 107476 182164 107528 182170
rect 107476 182106 107528 182112
rect 107660 182164 107712 182170
rect 107660 182106 107712 182112
rect 100666 173904 100722 173913
rect 100666 173839 100722 173848
rect 100850 173904 100906 173913
rect 100850 173839 100906 173848
rect 100864 164257 100892 173839
rect 107672 172553 107700 182106
rect 107474 172544 107530 172553
rect 107474 172479 107530 172488
rect 107658 172544 107714 172553
rect 107658 172479 107714 172488
rect 100666 164248 100722 164257
rect 100666 164183 100722 164192
rect 100850 164248 100906 164257
rect 100850 164183 100906 164192
rect 100680 154562 100708 164183
rect 107488 162858 107516 172479
rect 107476 162852 107528 162858
rect 107476 162794 107528 162800
rect 100668 154556 100720 154562
rect 100668 154498 100720 154504
rect 100852 154556 100904 154562
rect 100852 154498 100904 154504
rect 100864 144945 100892 154498
rect 107476 153264 107528 153270
rect 107476 153206 107528 153212
rect 100666 144936 100722 144945
rect 100666 144871 100722 144880
rect 100850 144936 100906 144945
rect 100850 144871 100906 144880
rect 100680 135250 100708 144871
rect 107488 143546 107516 153206
rect 107476 143540 107528 143546
rect 107476 143482 107528 143488
rect 100668 135244 100720 135250
rect 100668 135186 100720 135192
rect 100852 135244 100904 135250
rect 100852 135186 100904 135192
rect 100864 125633 100892 135186
rect 107476 133952 107528 133958
rect 107476 133894 107528 133900
rect 100666 125624 100722 125633
rect 100666 125559 100722 125568
rect 100850 125624 100906 125633
rect 100850 125559 100906 125568
rect 100680 115938 100708 125559
rect 107488 124166 107516 133894
rect 107476 124160 107528 124166
rect 107476 124102 107528 124108
rect 100668 115932 100720 115938
rect 100668 115874 100720 115880
rect 107476 114572 107528 114578
rect 107476 114514 107528 114520
rect 100668 106344 100720 106350
rect 100668 106286 100720 106292
rect 100680 96626 100708 106286
rect 107488 104854 107516 114514
rect 107476 104848 107528 104854
rect 107476 104790 107528 104796
rect 100668 96620 100720 96626
rect 100668 96562 100720 96568
rect 107476 95260 107528 95266
rect 107476 95202 107528 95208
rect 100668 87032 100720 87038
rect 100668 86974 100720 86980
rect 100680 77246 100708 86974
rect 107488 85542 107516 95202
rect 107476 85536 107528 85542
rect 107476 85478 107528 85484
rect 100668 77240 100720 77246
rect 100668 77182 100720 77188
rect 107476 75948 107528 75954
rect 107476 75890 107528 75896
rect 100668 67652 100720 67658
rect 100668 67594 100720 67600
rect 100680 57934 100708 67594
rect 107488 66230 107516 75890
rect 107476 66224 107528 66230
rect 107476 66166 107528 66172
rect 100668 57928 100720 57934
rect 100668 57870 100720 57876
rect 107476 56636 107528 56642
rect 107476 56578 107528 56584
rect 100668 48340 100720 48346
rect 100668 48282 100720 48288
rect 100680 38622 100708 48282
rect 107488 46918 107516 56578
rect 107476 46912 107528 46918
rect 107476 46854 107528 46860
rect 100668 38616 100720 38622
rect 100668 38558 100720 38564
rect 107476 37324 107528 37330
rect 107476 37266 107528 37272
rect 100668 29028 100720 29034
rect 100668 28970 100720 28976
rect 100680 19310 100708 28970
rect 107488 27606 107516 37266
rect 107476 27600 107528 27606
rect 107476 27542 107528 27548
rect 100484 19304 100536 19310
rect 100484 19246 100536 19252
rect 100668 19304 100720 19310
rect 100668 19246 100720 19252
rect 110328 19304 110380 19310
rect 110328 19246 110380 19252
rect 99288 19168 99340 19174
rect 99288 19110 99340 19116
rect 96528 19100 96580 19106
rect 96528 19042 96580 19048
rect 95148 15836 95200 15842
rect 95148 15778 95200 15784
rect 95160 3670 95188 15778
rect 96540 3670 96568 19042
rect 99196 15768 99248 15774
rect 99196 15710 99248 15716
rect 99208 3670 99236 15710
rect 93308 3664 93360 3670
rect 93308 3606 93360 3612
rect 93768 3664 93820 3670
rect 93768 3606 93820 3612
rect 94504 3664 94556 3670
rect 94504 3606 94556 3612
rect 95148 3664 95200 3670
rect 95148 3606 95200 3612
rect 95700 3664 95752 3670
rect 95700 3606 95752 3612
rect 96528 3664 96580 3670
rect 96528 3606 96580 3612
rect 98092 3664 98144 3670
rect 98092 3606 98144 3612
rect 99196 3664 99248 3670
rect 99196 3606 99248 3612
rect 92112 2848 92164 2854
rect 92112 2790 92164 2796
rect 92388 2848 92440 2854
rect 92388 2790 92440 2796
rect 90916 604 90968 610
rect 90916 546 90968 552
rect 90928 480 90956 546
rect 92124 480 92152 2790
rect 93320 480 93348 3606
rect 94516 480 94544 3606
rect 95712 480 95740 3606
rect 96896 3052 96948 3058
rect 96896 2994 96948 3000
rect 96908 480 96936 2994
rect 98104 480 98132 3606
rect 99300 480 99328 19110
rect 100496 9761 100524 19246
rect 103428 19236 103480 19242
rect 103428 19178 103480 19184
rect 102048 15700 102100 15706
rect 102048 15642 102100 15648
rect 100482 9752 100538 9761
rect 100482 9687 100538 9696
rect 100666 9752 100722 9761
rect 100666 9687 100722 9696
rect 100680 9654 100708 9687
rect 100668 9648 100720 9654
rect 100668 9590 100720 9596
rect 102060 3670 102088 15642
rect 103440 3670 103468 19178
rect 106188 15632 106240 15638
rect 106188 15574 106240 15580
rect 106200 3670 106228 15574
rect 108948 15564 109000 15570
rect 108948 15506 109000 15512
rect 107752 9716 107804 9722
rect 107752 9658 107804 9664
rect 106372 4752 106424 4758
rect 106372 4694 106424 4700
rect 101588 3664 101640 3670
rect 101588 3606 101640 3612
rect 102048 3664 102100 3670
rect 102048 3606 102100 3612
rect 102784 3664 102836 3670
rect 102784 3606 102836 3612
rect 103428 3664 103480 3670
rect 103428 3606 103480 3612
rect 105176 3664 105228 3670
rect 105176 3606 105228 3612
rect 106188 3664 106240 3670
rect 106188 3606 106240 3612
rect 100484 604 100536 610
rect 100484 546 100536 552
rect 100496 480 100524 546
rect 101600 480 101628 3606
rect 102796 480 102824 3606
rect 103980 3052 104032 3058
rect 103980 2994 104032 3000
rect 103992 480 104020 2994
rect 105188 480 105216 3606
rect 106384 480 106412 4694
rect 107764 610 107792 9658
rect 108960 9654 108988 15506
rect 108948 9648 109000 9654
rect 108948 9590 109000 9596
rect 110340 610 110368 19246
rect 113088 15496 113140 15502
rect 113088 15438 113140 15444
rect 113100 3670 113128 15438
rect 113548 5432 113600 5438
rect 113548 5374 113600 5380
rect 112352 3664 112404 3670
rect 112352 3606 112404 3612
rect 113088 3664 113140 3670
rect 113088 3606 113140 3612
rect 111156 2916 111208 2922
rect 111156 2858 111208 2864
rect 107568 604 107620 610
rect 107568 546 107620 552
rect 107752 604 107804 610
rect 107752 546 107804 552
rect 108764 604 108816 610
rect 108764 546 108816 552
rect 109960 604 110012 610
rect 109960 546 110012 552
rect 110328 604 110380 610
rect 110328 546 110380 552
rect 107580 480 107608 546
rect 108776 480 108804 546
rect 109972 480 110000 546
rect 111168 480 111196 2858
rect 112364 480 112392 3606
rect 113560 480 113588 5374
rect 115860 3670 115888 337146
rect 122748 337136 122800 337142
rect 122748 337078 122800 337084
rect 117228 15428 117280 15434
rect 117228 15370 117280 15376
rect 117240 3670 117268 15370
rect 119988 15360 120040 15366
rect 119988 15302 120040 15308
rect 120000 3670 120028 15302
rect 120632 4752 120684 4758
rect 120632 4694 120684 4700
rect 114744 3664 114796 3670
rect 114744 3606 114796 3612
rect 115848 3664 115900 3670
rect 115848 3606 115900 3612
rect 115940 3664 115992 3670
rect 115940 3606 115992 3612
rect 117228 3664 117280 3670
rect 117228 3606 117280 3612
rect 119436 3664 119488 3670
rect 119436 3606 119488 3612
rect 119988 3664 120040 3670
rect 119988 3606 120040 3612
rect 114756 480 114784 3606
rect 115952 480 115980 3606
rect 117136 2848 117188 2854
rect 117136 2790 117188 2796
rect 117148 480 117176 2790
rect 118240 2780 118292 2786
rect 118240 2722 118292 2728
rect 118252 480 118280 2722
rect 119448 480 119476 3606
rect 120644 480 120672 4694
rect 122760 3670 122788 337078
rect 173164 337068 173216 337074
rect 173164 337010 173216 337016
rect 124128 15292 124180 15298
rect 124128 15234 124180 15240
rect 124140 3670 124168 15234
rect 167092 9512 167144 9518
rect 167092 9454 167144 9460
rect 165896 9376 165948 9382
rect 165896 9318 165948 9324
rect 164700 9308 164752 9314
rect 164700 9250 164752 9256
rect 163504 9240 163556 9246
rect 163504 9182 163556 9188
rect 162308 9172 162360 9178
rect 162308 9114 162360 9120
rect 161112 9104 161164 9110
rect 161112 9046 161164 9052
rect 129004 9036 129056 9042
rect 129004 8978 129056 8984
rect 126612 8968 126664 8974
rect 126612 8910 126664 8916
rect 124220 5500 124272 5506
rect 124220 5442 124272 5448
rect 121828 3664 121880 3670
rect 121828 3606 121880 3612
rect 122748 3664 122800 3670
rect 122748 3606 122800 3612
rect 123024 3664 123076 3670
rect 123024 3606 123076 3612
rect 124128 3664 124180 3670
rect 124128 3606 124180 3612
rect 121840 480 121868 3606
rect 123036 480 123064 3606
rect 124232 480 124260 5442
rect 125416 5364 125468 5370
rect 125416 5306 125468 5312
rect 125428 480 125456 5306
rect 126624 480 126652 8910
rect 127808 4820 127860 4826
rect 127808 4762 127860 4768
rect 127820 480 127848 4762
rect 129016 480 129044 8978
rect 150438 8256 150494 8265
rect 150438 8191 150494 8200
rect 146850 8120 146906 8129
rect 146850 8055 146906 8064
rect 143262 7984 143318 7993
rect 143262 7919 143318 7928
rect 139674 7848 139730 7857
rect 139674 7783 139730 7792
rect 136086 7712 136142 7721
rect 136086 7647 136142 7656
rect 132590 7576 132646 7585
rect 132590 7511 132646 7520
rect 131394 6216 131450 6225
rect 131394 6151 131450 6160
rect 130198 4856 130254 4865
rect 130198 4791 130254 4800
rect 130212 480 130240 4791
rect 131408 480 131436 6151
rect 132604 480 132632 7511
rect 134890 6352 134946 6361
rect 134890 6287 134946 6296
rect 133788 4888 133840 4894
rect 133788 4830 133840 4836
rect 133800 480 133828 4830
rect 134904 480 134932 6287
rect 136100 480 136128 7647
rect 138478 6488 138534 6497
rect 138478 6423 138534 6432
rect 137282 4992 137338 5001
rect 137282 4927 137338 4936
rect 137296 480 137324 4927
rect 138492 480 138520 6423
rect 139688 480 139716 7783
rect 142066 6624 142122 6633
rect 142066 6559 142122 6568
rect 140872 4956 140924 4962
rect 140872 4898 140924 4904
rect 140884 480 140912 4898
rect 142080 480 142108 6559
rect 143276 480 143304 7919
rect 145654 6760 145710 6769
rect 145654 6695 145710 6704
rect 144460 5024 144512 5030
rect 144460 4966 144512 4972
rect 144472 480 144500 4966
rect 145668 480 145696 6695
rect 146864 480 146892 8055
rect 149242 6896 149298 6905
rect 149242 6831 149298 6840
rect 148048 5092 148100 5098
rect 148048 5034 148100 5040
rect 148060 480 148088 5034
rect 149256 480 149284 6831
rect 150452 480 150480 8191
rect 157524 7676 157576 7682
rect 157524 7618 157576 7624
rect 153936 7608 153988 7614
rect 153936 7550 153988 7556
rect 152740 6180 152792 6186
rect 152740 6122 152792 6128
rect 151544 5160 151596 5166
rect 151544 5102 151596 5108
rect 151556 480 151584 5102
rect 152752 480 152780 6122
rect 153948 480 153976 7550
rect 156328 6248 156380 6254
rect 156328 6190 156380 6196
rect 155132 5228 155184 5234
rect 155132 5170 155184 5176
rect 155144 480 155172 5170
rect 156340 480 156368 6190
rect 157536 480 157564 7618
rect 159916 6316 159968 6322
rect 159916 6258 159968 6264
rect 158720 5296 158772 5302
rect 158720 5238 158772 5244
rect 158732 480 158760 5238
rect 159928 480 159956 6258
rect 161124 480 161152 9046
rect 162320 480 162348 9114
rect 163516 480 163544 9182
rect 164712 480 164740 9250
rect 165908 480 165936 9318
rect 167104 480 167132 9454
rect 169392 9444 169444 9450
rect 169392 9386 169444 9392
rect 168196 7744 168248 7750
rect 168196 7686 168248 7692
rect 168208 480 168236 7686
rect 169404 480 169432 9386
rect 171784 7812 171836 7818
rect 171784 7754 171836 7760
rect 170588 6384 170640 6390
rect 170588 6326 170640 6332
rect 170600 480 170628 6326
rect 171796 480 171824 7754
rect 172980 4684 173032 4690
rect 172980 4626 173032 4632
rect 172992 480 173020 4626
rect 173176 4554 173204 337010
rect 182824 337000 182876 337006
rect 182824 336942 182876 336948
rect 182548 8016 182600 8022
rect 182548 7958 182600 7964
rect 178960 7948 179012 7954
rect 178960 7890 179012 7896
rect 175372 7880 175424 7886
rect 175372 7822 175424 7828
rect 174176 6452 174228 6458
rect 174176 6394 174228 6400
rect 173164 4548 173216 4554
rect 173164 4490 173216 4496
rect 174188 480 174216 6394
rect 175384 480 175412 7822
rect 177764 6520 177816 6526
rect 177764 6462 177816 6468
rect 176566 5128 176622 5137
rect 176566 5063 176622 5072
rect 176580 480 176608 5063
rect 177776 480 177804 6462
rect 178972 480 179000 7890
rect 181352 6588 181404 6594
rect 181352 6530 181404 6536
rect 180156 4616 180208 4622
rect 180156 4558 180208 4564
rect 180168 480 180196 4558
rect 180708 4344 180760 4350
rect 180708 4286 180760 4292
rect 180524 3868 180576 3874
rect 180524 3810 180576 3816
rect 180536 3754 180564 3810
rect 180536 3738 180656 3754
rect 180720 3738 180748 4286
rect 180536 3732 180668 3738
rect 180536 3726 180616 3732
rect 180616 3674 180668 3680
rect 180708 3732 180760 3738
rect 180708 3674 180760 3680
rect 181364 480 181392 6530
rect 182560 480 182588 7958
rect 182836 5438 182864 336942
rect 186964 336932 187016 336938
rect 186964 336874 187016 336880
rect 186044 8084 186096 8090
rect 186044 8026 186096 8032
rect 184848 6656 184900 6662
rect 184848 6598 184900 6604
rect 182824 5432 182876 5438
rect 182824 5374 182876 5380
rect 183742 5264 183798 5273
rect 183742 5199 183798 5208
rect 183756 480 183784 5199
rect 184860 480 184888 6598
rect 186056 480 186084 8026
rect 186976 4758 187004 336874
rect 191104 336864 191156 336870
rect 191104 336806 191156 336812
rect 189632 8152 189684 8158
rect 189632 8094 189684 8100
rect 188436 6724 188488 6730
rect 188436 6666 188488 6672
rect 187240 5432 187292 5438
rect 187240 5374 187292 5380
rect 186964 4752 187016 4758
rect 186964 4694 187016 4700
rect 187252 480 187280 5374
rect 188448 480 188476 6666
rect 189644 480 189672 8094
rect 191116 5506 191144 336806
rect 195244 336796 195296 336802
rect 195244 336738 195296 336744
rect 193220 8220 193272 8226
rect 193220 8162 193272 8168
rect 192024 6792 192076 6798
rect 192024 6734 192076 6740
rect 191104 5500 191156 5506
rect 191104 5442 191156 5448
rect 190826 5400 190882 5409
rect 190826 5335 190882 5344
rect 190840 480 190868 5335
rect 192036 480 192064 6734
rect 193232 480 193260 8162
rect 194416 5500 194468 5506
rect 194416 5442 194468 5448
rect 194428 480 194456 5442
rect 195256 5370 195284 336738
rect 229112 16833 229140 459326
rect 258814 459368 258870 459377
rect 234398 459326 234554 459354
rect 258750 459326 258814 459354
rect 234342 459303 234398 459312
rect 329012 459400 329064 459406
rect 324870 459368 324926 459377
rect 321704 459348 321954 459354
rect 321652 459342 321954 459348
rect 321664 459326 321954 459342
rect 258814 459303 258870 459312
rect 324926 459326 325082 459354
rect 325896 459338 326094 459354
rect 327920 459338 328210 459354
rect 345754 459368 345810 459377
rect 329064 459348 329314 459354
rect 329012 459342 329314 459348
rect 325884 459332 326094 459338
rect 324870 459303 324926 459312
rect 325936 459326 326094 459332
rect 327908 459332 328210 459338
rect 325884 459274 325936 459280
rect 327960 459326 328210 459332
rect 329024 459326 329314 459342
rect 331232 459338 331430 459354
rect 332152 459338 332442 459354
rect 334176 459338 334558 459354
rect 335372 459338 335570 459354
rect 337304 459338 337686 459354
rect 338408 459338 338790 459354
rect 340708 459338 340906 459354
rect 341536 459338 341918 459354
rect 331220 459332 331430 459338
rect 327908 459274 327960 459280
rect 331272 459326 331430 459332
rect 332140 459332 332442 459338
rect 331220 459274 331272 459280
rect 332192 459326 332442 459332
rect 334164 459332 334558 459338
rect 332140 459274 332192 459280
rect 334216 459326 334558 459332
rect 335360 459332 335570 459338
rect 334164 459274 334216 459280
rect 335412 459326 335570 459332
rect 337292 459332 337686 459338
rect 335360 459274 335412 459280
rect 337344 459326 337686 459332
rect 338396 459332 338790 459338
rect 337292 459274 337344 459280
rect 338448 459326 338790 459332
rect 340696 459332 340906 459338
rect 338396 459274 338448 459280
rect 340748 459326 340906 459332
rect 341524 459332 341918 459338
rect 340696 459274 340748 459280
rect 341576 459326 341918 459332
rect 347226 459368 347282 459377
rect 345810 459326 346150 459354
rect 347162 459326 347226 459354
rect 345754 459303 345810 459312
rect 349278 459326 349844 459354
rect 347226 459303 347282 459312
rect 341524 459274 341576 459280
rect 254242 340190 254440 340218
rect 262798 340190 262996 340218
rect 229296 340054 230046 340082
rect 230124 340054 230230 340082
rect 229192 335640 229244 335646
rect 229192 335582 229244 335588
rect 229098 16824 229154 16833
rect 229098 16759 229154 16768
rect 196808 8288 196860 8294
rect 196808 8230 196860 8236
rect 195612 6860 195664 6866
rect 195612 6802 195664 6808
rect 195244 5364 195296 5370
rect 195244 5306 195296 5312
rect 195624 480 195652 6802
rect 196820 480 196848 8230
rect 200396 7540 200448 7546
rect 200396 7482 200448 7488
rect 199200 6112 199252 6118
rect 199200 6054 199252 6060
rect 198004 5364 198056 5370
rect 198004 5306 198056 5312
rect 198016 480 198044 5306
rect 199212 480 199240 6054
rect 200408 480 200436 7482
rect 203892 7472 203944 7478
rect 203892 7414 203944 7420
rect 202696 6044 202748 6050
rect 202696 5986 202748 5992
rect 201500 4752 201552 4758
rect 201500 4694 201552 4700
rect 201512 480 201540 4694
rect 202708 480 202736 5986
rect 203904 480 203932 7414
rect 207480 7404 207532 7410
rect 207480 7346 207532 7352
rect 206284 5976 206336 5982
rect 206284 5918 206336 5924
rect 205086 5536 205142 5545
rect 205086 5471 205142 5480
rect 205100 480 205128 5471
rect 206296 480 206324 5918
rect 207492 480 207520 7346
rect 211068 7336 211120 7342
rect 211068 7278 211120 7284
rect 209872 5908 209924 5914
rect 209872 5850 209924 5856
rect 208676 4548 208728 4554
rect 208676 4490 208728 4496
rect 208688 480 208716 4490
rect 209884 480 209912 5850
rect 211080 480 211108 7278
rect 214656 7268 214708 7274
rect 214656 7210 214708 7216
rect 213460 5840 213512 5846
rect 213460 5782 213512 5788
rect 212264 4480 212316 4486
rect 212264 4422 212316 4428
rect 212276 480 212304 4422
rect 213472 480 213500 5782
rect 214668 480 214696 7210
rect 218152 7200 218204 7206
rect 218152 7142 218204 7148
rect 217048 5772 217100 5778
rect 217048 5714 217100 5720
rect 215852 4412 215904 4418
rect 215852 4354 215904 4360
rect 215864 480 215892 4354
rect 217060 480 217088 5714
rect 218164 480 218192 7142
rect 221740 7132 221792 7138
rect 221740 7074 221792 7080
rect 220544 5704 220596 5710
rect 220544 5646 220596 5652
rect 219348 4344 219400 4350
rect 219348 4286 219400 4292
rect 219360 480 219388 4286
rect 220556 480 220584 5646
rect 221752 480 221780 7074
rect 225328 7064 225380 7070
rect 225328 7006 225380 7012
rect 224132 5636 224184 5642
rect 224132 5578 224184 5584
rect 222936 4276 222988 4282
rect 222936 4218 222988 4224
rect 222948 480 222976 4218
rect 224144 480 224172 5578
rect 224776 3664 224828 3670
rect 224776 3606 224828 3612
rect 224960 3664 225012 3670
rect 224960 3606 225012 3612
rect 224788 3233 224816 3606
rect 224972 3233 225000 3606
rect 224774 3224 224830 3233
rect 224774 3159 224830 3168
rect 224958 3224 225014 3233
rect 224958 3159 225014 3168
rect 225340 480 225368 7006
rect 228916 6996 228968 7002
rect 228916 6938 228968 6944
rect 227720 5568 227772 5574
rect 227720 5510 227772 5516
rect 226524 4208 226576 4214
rect 226524 4150 226576 4156
rect 226536 480 226564 4150
rect 227732 480 227760 5510
rect 228928 480 228956 6938
rect 229204 4826 229232 335582
rect 229296 8974 229324 340054
rect 230124 335646 230152 340054
rect 230112 335640 230164 335646
rect 230112 335582 230164 335588
rect 230492 9042 230520 340068
rect 230584 340054 230690 340082
rect 230768 340054 230966 340082
rect 231044 340054 231242 340082
rect 231320 340054 231426 340082
rect 231596 340054 231702 340082
rect 230480 9036 230532 9042
rect 230480 8978 230532 8984
rect 229284 8968 229336 8974
rect 229284 8910 229336 8916
rect 230584 4865 230612 340054
rect 230768 6225 230796 340054
rect 231044 335730 231072 340054
rect 231214 338056 231270 338065
rect 231214 337991 231270 338000
rect 230860 335702 231072 335730
rect 230860 7585 230888 335702
rect 231032 331900 231084 331906
rect 231032 331842 231084 331848
rect 230846 7576 230902 7585
rect 230846 7511 230902 7520
rect 230754 6216 230810 6225
rect 230754 6151 230810 6160
rect 231044 4894 231072 331842
rect 231228 328522 231256 337991
rect 231320 331906 231348 340054
rect 231596 338065 231624 340054
rect 231860 338700 231912 338706
rect 231860 338642 231912 338648
rect 231582 338056 231638 338065
rect 231582 337991 231638 338000
rect 231308 331900 231360 331906
rect 231308 331842 231360 331848
rect 231136 328494 231256 328522
rect 231136 328438 231164 328494
rect 231124 328432 231176 328438
rect 231124 328374 231176 328380
rect 231216 318844 231268 318850
rect 231216 318786 231268 318792
rect 231228 311982 231256 318786
rect 231216 311976 231268 311982
rect 231216 311918 231268 311924
rect 231216 311772 231268 311778
rect 231216 311714 231268 311720
rect 231228 299470 231256 311714
rect 231216 299464 231268 299470
rect 231216 299406 231268 299412
rect 231216 289876 231268 289882
rect 231216 289818 231268 289824
rect 231228 280158 231256 289818
rect 231216 280152 231268 280158
rect 231216 280094 231268 280100
rect 231216 270564 231268 270570
rect 231216 270506 231268 270512
rect 231228 260846 231256 270506
rect 231768 262948 231820 262954
rect 231768 262890 231820 262896
rect 231216 260840 231268 260846
rect 231216 260782 231268 260788
rect 231780 258097 231808 262890
rect 231766 258088 231822 258097
rect 231766 258023 231822 258032
rect 231216 251252 231268 251258
rect 231216 251194 231268 251200
rect 231228 241505 231256 251194
rect 231214 241496 231270 241505
rect 231214 241431 231270 241440
rect 231398 241496 231454 241505
rect 231398 241431 231454 241440
rect 231412 231878 231440 241431
rect 231216 231872 231268 231878
rect 231216 231814 231268 231820
rect 231400 231872 231452 231878
rect 231400 231814 231452 231820
rect 231228 222193 231256 231814
rect 231214 222184 231270 222193
rect 231214 222119 231270 222128
rect 231398 222184 231454 222193
rect 231398 222119 231454 222128
rect 231412 212566 231440 222119
rect 231216 212560 231268 212566
rect 231216 212502 231268 212508
rect 231400 212560 231452 212566
rect 231400 212502 231452 212508
rect 231228 202881 231256 212502
rect 231214 202872 231270 202881
rect 231214 202807 231270 202816
rect 231398 202872 231454 202881
rect 231398 202807 231454 202816
rect 231412 193254 231440 202807
rect 231216 193248 231268 193254
rect 231216 193190 231268 193196
rect 231400 193248 231452 193254
rect 231400 193190 231452 193196
rect 231228 183569 231256 193190
rect 231214 183560 231270 183569
rect 231214 183495 231270 183504
rect 231398 183560 231454 183569
rect 231398 183495 231454 183504
rect 231412 173942 231440 183495
rect 231216 173936 231268 173942
rect 231216 173878 231268 173884
rect 231400 173936 231452 173942
rect 231400 173878 231452 173884
rect 231228 157350 231256 173878
rect 231216 157344 231268 157350
rect 231216 157286 231268 157292
rect 231216 157208 231268 157214
rect 231216 157150 231268 157156
rect 231228 154562 231256 157150
rect 231216 154556 231268 154562
rect 231216 154498 231268 154504
rect 231400 154556 231452 154562
rect 231400 154498 231452 154504
rect 231412 144945 231440 154498
rect 231214 144936 231270 144945
rect 231214 144871 231270 144880
rect 231398 144936 231454 144945
rect 231398 144871 231454 144880
rect 231228 138038 231256 144871
rect 231216 138032 231268 138038
rect 231216 137974 231268 137980
rect 231216 135380 231268 135386
rect 231216 135322 231268 135328
rect 231228 135250 231256 135322
rect 231216 135244 231268 135250
rect 231216 135186 231268 135192
rect 231400 135244 231452 135250
rect 231400 135186 231452 135192
rect 231412 125633 231440 135186
rect 231214 125624 231270 125633
rect 231214 125559 231270 125568
rect 231398 125624 231454 125633
rect 231398 125559 231454 125568
rect 231228 118726 231256 125559
rect 231216 118720 231268 118726
rect 231216 118662 231268 118668
rect 231216 116068 231268 116074
rect 231216 116010 231268 116016
rect 231228 115938 231256 116010
rect 231216 115932 231268 115938
rect 231216 115874 231268 115880
rect 231216 106344 231268 106350
rect 231216 106286 231268 106292
rect 231228 99414 231256 106286
rect 231216 99408 231268 99414
rect 231216 99350 231268 99356
rect 231216 96756 231268 96762
rect 231216 96698 231268 96704
rect 231228 80170 231256 96698
rect 231216 80164 231268 80170
rect 231216 80106 231268 80112
rect 231216 80028 231268 80034
rect 231216 79970 231268 79976
rect 231228 70394 231256 79970
rect 231228 70366 231348 70394
rect 231320 67658 231348 70366
rect 231124 67652 231176 67658
rect 231124 67594 231176 67600
rect 231308 67652 231360 67658
rect 231308 67594 231360 67600
rect 231136 66230 231164 67594
rect 231124 66224 231176 66230
rect 231124 66166 231176 66172
rect 231308 66224 231360 66230
rect 231308 66166 231360 66172
rect 231320 55214 231348 66166
rect 231308 55208 231360 55214
rect 231308 55150 231360 55156
rect 231308 45620 231360 45626
rect 231308 45562 231360 45568
rect 231320 40746 231348 45562
rect 231228 40718 231348 40746
rect 231228 32450 231256 40718
rect 231136 32422 231256 32450
rect 231136 16674 231164 32422
rect 231136 16646 231256 16674
rect 231228 12594 231256 16646
rect 231228 12566 231348 12594
rect 231320 9228 231348 12566
rect 231228 9200 231348 9228
rect 231228 6361 231256 9200
rect 231214 6352 231270 6361
rect 231214 6287 231270 6296
rect 231872 5001 231900 338642
rect 231964 335646 231992 340068
rect 232148 338706 232176 340068
rect 232240 340054 232438 340082
rect 232516 340054 232714 340082
rect 232792 340054 232898 340082
rect 232136 338700 232188 338706
rect 232136 338642 232188 338648
rect 232240 335782 232268 340054
rect 232228 335776 232280 335782
rect 232228 335718 232280 335724
rect 232516 335696 232544 340054
rect 232424 335668 232544 335696
rect 231952 335640 232004 335646
rect 231952 335582 232004 335588
rect 232228 335640 232280 335646
rect 232228 335582 232280 335588
rect 232136 328500 232188 328506
rect 232136 328442 232188 328448
rect 232148 318866 232176 328442
rect 232056 318838 232176 318866
rect 232056 311964 232084 318838
rect 231964 311936 232084 311964
rect 231964 311794 231992 311936
rect 231964 311766 232084 311794
rect 232056 299470 232084 311766
rect 231952 299464 232004 299470
rect 231952 299406 232004 299412
rect 232044 299464 232096 299470
rect 232044 299406 232096 299412
rect 231964 298110 231992 299406
rect 231952 298104 232004 298110
rect 231952 298046 232004 298052
rect 232044 298104 232096 298110
rect 232044 298046 232096 298052
rect 232056 280158 232084 298046
rect 232044 280152 232096 280158
rect 232044 280094 232096 280100
rect 232136 280152 232188 280158
rect 232136 280094 232188 280100
rect 232148 278769 232176 280094
rect 231950 278760 232006 278769
rect 231950 278695 232006 278704
rect 232134 278760 232190 278769
rect 232134 278695 232190 278704
rect 231964 269142 231992 278695
rect 231952 269136 232004 269142
rect 231952 269078 232004 269084
rect 232136 269136 232188 269142
rect 232136 269078 232188 269084
rect 232148 267730 232176 269078
rect 232056 267702 232176 267730
rect 232056 262954 232084 267702
rect 232044 262948 232096 262954
rect 232044 262890 232096 262896
rect 231950 258088 232006 258097
rect 232006 258058 232084 258074
rect 232006 258052 232096 258058
rect 232006 258046 232044 258052
rect 231950 258023 232006 258032
rect 232044 257994 232096 258000
rect 232136 253904 232188 253910
rect 232136 253846 232188 253852
rect 232148 240174 232176 253846
rect 232044 240168 232096 240174
rect 232044 240110 232096 240116
rect 232136 240168 232188 240174
rect 232136 240110 232188 240116
rect 232056 234666 232084 240110
rect 232044 234660 232096 234666
rect 232044 234602 232096 234608
rect 232044 230512 232096 230518
rect 232044 230454 232096 230460
rect 232056 225010 232084 230454
rect 232044 225004 232096 225010
rect 232044 224946 232096 224952
rect 232044 222216 232096 222222
rect 232044 222158 232096 222164
rect 232056 220833 232084 222158
rect 232042 220824 232098 220833
rect 232042 220759 232098 220768
rect 232042 211168 232098 211177
rect 232042 211103 232098 211112
rect 232056 202881 232084 211103
rect 232042 202872 232098 202881
rect 232042 202807 232098 202816
rect 232134 202736 232190 202745
rect 232134 202671 232190 202680
rect 232148 197962 232176 202671
rect 232056 197934 232176 197962
rect 232056 182170 232084 197934
rect 232136 191820 232188 191826
rect 232136 191762 232188 191768
rect 232148 182209 232176 191762
rect 232134 182200 232190 182209
rect 232044 182164 232096 182170
rect 232134 182135 232190 182144
rect 232044 182106 232096 182112
rect 231952 182096 232004 182102
rect 231952 182038 232004 182044
rect 231964 172553 231992 182038
rect 231950 172544 232006 172553
rect 231950 172479 232006 172488
rect 232134 172544 232190 172553
rect 232134 172479 232190 172488
rect 232148 167686 232176 172479
rect 231952 167680 232004 167686
rect 231952 167622 232004 167628
rect 232136 167680 232188 167686
rect 232136 167622 232188 167628
rect 231964 166818 231992 167622
rect 231964 166790 232084 166818
rect 232056 162858 232084 166790
rect 232044 162852 232096 162858
rect 232044 162794 232096 162800
rect 232136 162852 232188 162858
rect 232136 162794 232188 162800
rect 232148 153202 232176 162794
rect 232136 153196 232188 153202
rect 232136 153138 232188 153144
rect 232044 143608 232096 143614
rect 232044 143550 232096 143556
rect 232056 142118 232084 143550
rect 232044 142112 232096 142118
rect 232044 142054 232096 142060
rect 232136 132524 232188 132530
rect 232136 132466 232188 132472
rect 232148 111790 232176 132466
rect 232044 111784 232096 111790
rect 232044 111726 232096 111732
rect 232136 111784 232188 111790
rect 232136 111726 232188 111732
rect 232056 103476 232084 111726
rect 232056 103448 232176 103476
rect 232148 102134 232176 103448
rect 232136 102128 232188 102134
rect 232136 102070 232188 102076
rect 232136 92540 232188 92546
rect 232136 92482 232188 92488
rect 232148 81462 232176 92482
rect 232240 85406 232268 335582
rect 232424 328522 232452 335668
rect 232792 335594 232820 340054
rect 233160 338842 233188 340068
rect 232872 338836 232924 338842
rect 232872 338778 232924 338784
rect 233148 338836 233200 338842
rect 233148 338778 233200 338784
rect 232332 328494 232452 328522
rect 232516 335566 232820 335594
rect 232332 318850 232360 328494
rect 232320 318844 232372 318850
rect 232320 318786 232372 318792
rect 232412 318844 232464 318850
rect 232412 318786 232464 318792
rect 232424 317422 232452 318786
rect 232320 317416 232372 317422
rect 232320 317358 232372 317364
rect 232412 317416 232464 317422
rect 232412 317358 232464 317364
rect 232332 299470 232360 317358
rect 232320 299464 232372 299470
rect 232320 299406 232372 299412
rect 232412 299464 232464 299470
rect 232412 299406 232464 299412
rect 232424 298110 232452 299406
rect 232412 298104 232464 298110
rect 232412 298046 232464 298052
rect 232412 288448 232464 288454
rect 232412 288390 232464 288396
rect 232424 260930 232452 288390
rect 232332 260902 232452 260930
rect 232332 258058 232360 260902
rect 232320 258052 232372 258058
rect 232320 257994 232372 258000
rect 232320 253224 232372 253230
rect 232320 253166 232372 253172
rect 232332 240145 232360 253166
rect 232318 240136 232374 240145
rect 232318 240071 232374 240080
rect 232320 222284 232372 222290
rect 232320 222226 232372 222232
rect 232332 220833 232360 222226
rect 232318 220824 232374 220833
rect 232318 220759 232374 220768
rect 232320 202904 232372 202910
rect 232320 202846 232372 202852
rect 232332 193254 232360 202846
rect 232320 193248 232372 193254
rect 232320 193190 232372 193196
rect 232412 193248 232464 193254
rect 232412 193190 232464 193196
rect 232424 191826 232452 193190
rect 232412 191820 232464 191826
rect 232412 191762 232464 191768
rect 232318 182200 232374 182209
rect 232318 182135 232320 182144
rect 232372 182135 232374 182144
rect 232320 182106 232372 182112
rect 232412 172576 232464 172582
rect 232412 172518 232464 172524
rect 232424 167074 232452 172518
rect 232412 167068 232464 167074
rect 232412 167010 232464 167016
rect 232320 167000 232372 167006
rect 232320 166942 232372 166948
rect 232332 162858 232360 166942
rect 232320 162852 232372 162858
rect 232320 162794 232372 162800
rect 232516 139641 232544 335566
rect 232884 333282 232912 338778
rect 233332 335708 233384 335714
rect 233332 335650 233384 335656
rect 233240 335640 233292 335646
rect 233240 335582 233292 335588
rect 232608 333254 232912 333282
rect 232608 318850 232636 333254
rect 232596 318844 232648 318850
rect 232596 318786 232648 318792
rect 232688 318844 232740 318850
rect 232688 318786 232740 318792
rect 232700 292670 232728 318786
rect 232688 292664 232740 292670
rect 232688 292606 232740 292612
rect 232688 292528 232740 292534
rect 232688 292470 232740 292476
rect 232700 273358 232728 292470
rect 232688 273352 232740 273358
rect 232688 273294 232740 273300
rect 232688 273216 232740 273222
rect 232688 273158 232740 273164
rect 232700 253994 232728 273158
rect 232608 253966 232728 253994
rect 232608 253858 232636 253966
rect 232608 253830 232728 253858
rect 232594 240136 232650 240145
rect 232700 240106 232728 253830
rect 232594 240071 232650 240080
rect 232688 240100 232740 240106
rect 232608 222290 232636 240071
rect 232688 240042 232740 240048
rect 232688 235340 232740 235346
rect 232688 235282 232740 235288
rect 232596 222284 232648 222290
rect 232596 222226 232648 222232
rect 232700 215370 232728 235282
rect 232778 220824 232834 220833
rect 232778 220759 232834 220768
rect 232608 215342 232728 215370
rect 232608 215234 232636 215342
rect 232608 215206 232728 215234
rect 232596 215144 232648 215150
rect 232596 215086 232648 215092
rect 232608 202910 232636 215086
rect 232596 202904 232648 202910
rect 232596 202846 232648 202852
rect 232700 202858 232728 215206
rect 232792 215150 232820 220759
rect 232780 215144 232832 215150
rect 232780 215086 232832 215092
rect 232700 202830 232820 202858
rect 232792 196042 232820 202830
rect 232780 196036 232832 196042
rect 232780 195978 232832 195984
rect 232688 195968 232740 195974
rect 232688 195910 232740 195916
rect 232700 176662 232728 195910
rect 232688 176656 232740 176662
rect 232688 176598 232740 176604
rect 232688 176520 232740 176526
rect 232688 176462 232740 176468
rect 232596 162852 232648 162858
rect 232596 162794 232648 162800
rect 232608 161430 232636 162794
rect 232596 161424 232648 161430
rect 232596 161366 232648 161372
rect 232596 153196 232648 153202
rect 232596 153138 232648 153144
rect 232502 139632 232558 139641
rect 232502 139567 232558 139576
rect 232502 139496 232558 139505
rect 232502 139431 232558 139440
rect 232412 139392 232464 139398
rect 232412 139334 232464 139340
rect 232424 136610 232452 139334
rect 232412 136604 232464 136610
rect 232412 136546 232464 136552
rect 232412 118720 232464 118726
rect 232412 118662 232464 118668
rect 232424 113098 232452 118662
rect 232332 113070 232452 113098
rect 232332 107030 232360 113070
rect 232320 107024 232372 107030
rect 232320 106966 232372 106972
rect 232320 93900 232372 93906
rect 232320 93842 232372 93848
rect 232332 89758 232360 93842
rect 232320 89752 232372 89758
rect 232320 89694 232372 89700
rect 232228 85400 232280 85406
rect 232228 85342 232280 85348
rect 232228 85264 232280 85270
rect 232228 85206 232280 85212
rect 232044 81456 232096 81462
rect 232044 81398 232096 81404
rect 232136 81456 232188 81462
rect 232136 81398 232188 81404
rect 232056 73114 232084 81398
rect 232056 73098 232176 73114
rect 232056 73092 232188 73098
rect 232056 73086 232136 73092
rect 232136 73034 232188 73040
rect 232136 46980 232188 46986
rect 232136 46922 232188 46928
rect 232148 19258 232176 46922
rect 232056 19230 232176 19258
rect 232056 6497 232084 19230
rect 232240 7721 232268 85206
rect 232412 75948 232464 75954
rect 232412 75890 232464 75896
rect 232424 67674 232452 75890
rect 232332 67646 232452 67674
rect 232332 66230 232360 67646
rect 232320 66224 232372 66230
rect 232320 66166 232372 66172
rect 232412 66224 232464 66230
rect 232412 66166 232464 66172
rect 232424 40730 232452 66166
rect 232412 40724 232464 40730
rect 232412 40666 232464 40672
rect 232320 27668 232372 27674
rect 232320 27610 232372 27616
rect 232332 7857 232360 27610
rect 232318 7848 232374 7857
rect 232318 7783 232374 7792
rect 232226 7712 232282 7721
rect 232226 7647 232282 7656
rect 232042 6488 232098 6497
rect 232042 6423 232098 6432
rect 232516 5080 232544 139431
rect 232608 139398 232636 153138
rect 232596 139392 232648 139398
rect 232596 139334 232648 139340
rect 232700 138106 232728 176462
rect 232596 138100 232648 138106
rect 232596 138042 232648 138048
rect 232688 138100 232740 138106
rect 232688 138042 232740 138048
rect 232608 136649 232636 138042
rect 232594 136640 232650 136649
rect 232594 136575 232650 136584
rect 232870 136640 232926 136649
rect 232870 136575 232926 136584
rect 232884 127090 232912 136575
rect 232872 127084 232924 127090
rect 232872 127026 232924 127032
rect 232688 127016 232740 127022
rect 232688 126958 232740 126964
rect 232608 118726 232636 118757
rect 232700 118726 232728 126958
rect 232596 118720 232648 118726
rect 232688 118720 232740 118726
rect 232648 118668 232688 118674
rect 232596 118662 232740 118668
rect 232608 118646 232728 118662
rect 232700 117298 232728 118646
rect 232688 117292 232740 117298
rect 232688 117234 232740 117240
rect 232872 117224 232924 117230
rect 232872 117166 232924 117172
rect 232884 107681 232912 117166
rect 232686 107672 232742 107681
rect 232686 107607 232742 107616
rect 232870 107672 232926 107681
rect 232870 107607 232926 107616
rect 232700 99482 232728 107607
rect 232688 99476 232740 99482
rect 232688 99418 232740 99424
rect 232688 99340 232740 99346
rect 232688 99282 232740 99288
rect 232700 67658 232728 99282
rect 232596 67652 232648 67658
rect 232596 67594 232648 67600
rect 232688 67652 232740 67658
rect 232688 67594 232740 67600
rect 232608 51762 232636 67594
rect 232608 51734 232820 51762
rect 232792 40730 232820 51734
rect 232780 40724 232832 40730
rect 232780 40666 232832 40672
rect 232780 27668 232832 27674
rect 232780 27610 232832 27616
rect 232792 9722 232820 27610
rect 232596 9716 232648 9722
rect 232596 9658 232648 9664
rect 232780 9716 232832 9722
rect 232780 9658 232832 9664
rect 232608 6633 232636 9658
rect 232594 6624 232650 6633
rect 232594 6559 232650 6568
rect 232424 5052 232544 5080
rect 231858 4992 231914 5001
rect 232424 4962 232452 5052
rect 233252 5030 233280 335582
rect 233344 5098 233372 335650
rect 233436 7993 233464 340068
rect 233528 340054 233634 340082
rect 233712 340054 233910 340082
rect 233988 340054 234186 340082
rect 234264 340054 234370 340082
rect 234646 340054 234844 340082
rect 233528 335646 233556 340054
rect 233516 335640 233568 335646
rect 233516 335582 233568 335588
rect 233516 335504 233568 335510
rect 233516 335446 233568 335452
rect 233528 8129 233556 335446
rect 233514 8120 233570 8129
rect 233514 8055 233570 8064
rect 233422 7984 233478 7993
rect 233422 7919 233478 7928
rect 233712 6769 233740 340054
rect 233988 335510 234016 340054
rect 234264 335714 234292 340054
rect 234252 335708 234304 335714
rect 234252 335650 234304 335656
rect 234712 335640 234764 335646
rect 234712 335582 234764 335588
rect 233976 335504 234028 335510
rect 233976 335446 234028 335452
rect 233698 6760 233754 6769
rect 233698 6695 233754 6704
rect 234724 5166 234752 335582
rect 234816 6905 234844 340054
rect 234908 8265 234936 340068
rect 235000 340054 235106 340082
rect 235276 340054 235382 340082
rect 235460 340054 235658 340082
rect 235736 340054 235842 340082
rect 235000 335646 235028 340054
rect 234988 335640 235040 335646
rect 234988 335582 235040 335588
rect 235172 335640 235224 335646
rect 235172 335582 235224 335588
rect 234988 335504 235040 335510
rect 234988 335446 235040 335452
rect 234894 8256 234950 8265
rect 234894 8191 234950 8200
rect 235000 7614 235028 335446
rect 234988 7608 235040 7614
rect 234988 7550 235040 7556
rect 234802 6896 234858 6905
rect 234802 6831 234858 6840
rect 235184 5234 235212 335582
rect 235276 6186 235304 340054
rect 235460 335510 235488 340054
rect 235736 335646 235764 340054
rect 236000 335912 236052 335918
rect 236000 335854 236052 335860
rect 235724 335640 235776 335646
rect 235724 335582 235776 335588
rect 235448 335504 235500 335510
rect 235448 335446 235500 335452
rect 235264 6180 235316 6186
rect 235264 6122 235316 6128
rect 236012 5386 236040 335854
rect 236104 6254 236132 340068
rect 236288 340054 236394 340082
rect 236472 340054 236578 340082
rect 236656 340054 236854 340082
rect 236932 340054 237130 340082
rect 237208 340054 237314 340082
rect 237590 340054 237696 340082
rect 236184 335844 236236 335850
rect 236184 335786 236236 335792
rect 236196 6322 236224 335786
rect 236288 7682 236316 340054
rect 236472 335918 236500 340054
rect 236460 335912 236512 335918
rect 236460 335854 236512 335860
rect 236656 335850 236684 340054
rect 236644 335844 236696 335850
rect 236644 335786 236696 335792
rect 236932 335696 236960 340054
rect 236472 335668 236960 335696
rect 236472 9110 236500 335668
rect 237208 332722 237236 340054
rect 237380 335708 237432 335714
rect 237380 335650 237432 335656
rect 236736 332716 236788 332722
rect 236736 332658 236788 332664
rect 237196 332716 237248 332722
rect 237196 332658 237248 332664
rect 236748 24154 236776 332658
rect 236656 24126 236776 24154
rect 236656 9178 236684 24126
rect 236644 9172 236696 9178
rect 236644 9114 236696 9120
rect 236460 9104 236512 9110
rect 236460 9046 236512 9052
rect 237392 7750 237420 335650
rect 237472 335640 237524 335646
rect 237472 335582 237524 335588
rect 237484 9382 237512 335582
rect 237472 9376 237524 9382
rect 237472 9318 237524 9324
rect 237668 9246 237696 340054
rect 237760 340054 237866 340082
rect 237944 340054 238050 340082
rect 237760 9314 237788 340054
rect 237944 335646 237972 340054
rect 238312 338706 238340 340068
rect 238404 340054 238602 340082
rect 238786 340054 238892 340082
rect 238024 338700 238076 338706
rect 238024 338642 238076 338648
rect 238300 338700 238352 338706
rect 238300 338642 238352 338648
rect 237932 335640 237984 335646
rect 237932 335582 237984 335588
rect 238036 309126 238064 338642
rect 238404 335714 238432 340054
rect 238392 335708 238444 335714
rect 238392 335650 238444 335656
rect 238864 335442 238892 340054
rect 238956 340054 239062 340082
rect 238852 335436 238904 335442
rect 238852 335378 238904 335384
rect 238852 335300 238904 335306
rect 238852 335242 238904 335248
rect 238024 309120 238076 309126
rect 238024 309062 238076 309068
rect 238024 299532 238076 299538
rect 238024 299474 238076 299480
rect 238036 289814 238064 299474
rect 238024 289808 238076 289814
rect 238024 289750 238076 289756
rect 238024 280220 238076 280226
rect 238024 280162 238076 280168
rect 238036 270502 238064 280162
rect 238024 270496 238076 270502
rect 238024 270438 238076 270444
rect 238024 260908 238076 260914
rect 238024 260850 238076 260856
rect 238036 240145 238064 260850
rect 237838 240136 237894 240145
rect 237838 240071 237894 240080
rect 238022 240136 238078 240145
rect 238022 240071 238078 240080
rect 237852 230518 237880 240071
rect 237840 230512 237892 230518
rect 237840 230454 237892 230460
rect 237932 230512 237984 230518
rect 237932 230454 237984 230460
rect 237944 222222 237972 230454
rect 237932 222216 237984 222222
rect 237932 222158 237984 222164
rect 238024 222216 238076 222222
rect 238024 222158 238076 222164
rect 238036 212514 238064 222158
rect 238036 212486 238156 212514
rect 238128 202910 238156 212486
rect 238024 202904 238076 202910
rect 238024 202846 238076 202852
rect 238116 202904 238168 202910
rect 238116 202846 238168 202852
rect 238036 193202 238064 202846
rect 238036 193174 238156 193202
rect 238128 183598 238156 193174
rect 238024 183592 238076 183598
rect 238024 183534 238076 183540
rect 238116 183592 238168 183598
rect 238116 183534 238168 183540
rect 238036 19378 238064 183534
rect 238666 90536 238722 90545
rect 238666 90471 238722 90480
rect 238680 87145 238708 90471
rect 238666 87136 238722 87145
rect 238666 87071 238722 87080
rect 237932 19372 237984 19378
rect 237932 19314 237984 19320
rect 238024 19372 238076 19378
rect 238024 19314 238076 19320
rect 237944 9518 237972 19314
rect 237932 9512 237984 9518
rect 237932 9454 237984 9460
rect 237748 9308 237800 9314
rect 237748 9250 237800 9256
rect 237656 9240 237708 9246
rect 237656 9182 237708 9188
rect 237380 7744 237432 7750
rect 237380 7686 237432 7692
rect 236276 7676 236328 7682
rect 236276 7618 236328 7624
rect 238864 6458 238892 335242
rect 238852 6452 238904 6458
rect 238852 6394 238904 6400
rect 238956 6390 238984 340054
rect 239128 335640 239180 335646
rect 239128 335582 239180 335588
rect 239140 7886 239168 335582
rect 239220 335436 239272 335442
rect 239220 335378 239272 335384
rect 239232 9450 239260 335378
rect 239220 9444 239272 9450
rect 239220 9386 239272 9392
rect 239128 7880 239180 7886
rect 239128 7822 239180 7828
rect 239324 7818 239352 340068
rect 239416 340054 239522 340082
rect 239600 340054 239798 340082
rect 239876 340054 240074 340082
rect 240152 340054 240258 340082
rect 240336 340054 240534 340082
rect 239312 7812 239364 7818
rect 239312 7754 239364 7760
rect 238944 6384 238996 6390
rect 238944 6326 238996 6332
rect 236184 6316 236236 6322
rect 236184 6258 236236 6264
rect 236092 6248 236144 6254
rect 236092 6190 236144 6196
rect 235920 5358 236040 5386
rect 235920 5302 235948 5358
rect 235908 5296 235960 5302
rect 235908 5238 235960 5244
rect 236000 5296 236052 5302
rect 236000 5238 236052 5244
rect 235172 5228 235224 5234
rect 235172 5170 235224 5176
rect 234712 5160 234764 5166
rect 234712 5102 234764 5108
rect 233332 5092 233384 5098
rect 233332 5034 233384 5040
rect 234804 5092 234856 5098
rect 234804 5034 234856 5040
rect 233240 5024 233292 5030
rect 233240 4966 233292 4972
rect 233700 5024 233752 5030
rect 233700 4966 233752 4972
rect 231858 4927 231914 4936
rect 232412 4956 232464 4962
rect 232412 4898 232464 4904
rect 232504 4956 232556 4962
rect 232504 4898 232556 4904
rect 231032 4888 231084 4894
rect 230570 4856 230626 4865
rect 229192 4820 229244 4826
rect 229192 4762 229244 4768
rect 230112 4820 230164 4826
rect 231032 4830 231084 4836
rect 231308 4888 231360 4894
rect 231308 4830 231360 4836
rect 230570 4791 230626 4800
rect 230112 4762 230164 4768
rect 230124 480 230152 4762
rect 231320 480 231348 4830
rect 232516 480 232544 4898
rect 233712 480 233740 4966
rect 234816 480 234844 5034
rect 236012 480 236040 5238
rect 238392 5228 238444 5234
rect 238392 5170 238444 5176
rect 237196 5160 237248 5166
rect 237196 5102 237248 5108
rect 237208 480 237236 5102
rect 238404 480 238432 5170
rect 239416 4690 239444 340054
rect 239600 335306 239628 340054
rect 239876 335646 239904 340054
rect 239864 335640 239916 335646
rect 239864 335582 239916 335588
rect 239588 335300 239640 335306
rect 239588 335242 239640 335248
rect 240152 5137 240180 340054
rect 240232 37256 240284 37262
rect 240232 37198 240284 37204
rect 240244 18018 240272 37198
rect 240232 18012 240284 18018
rect 240232 17954 240284 17960
rect 240336 6526 240364 340054
rect 240416 335640 240468 335646
rect 240416 335582 240468 335588
rect 240428 6594 240456 335582
rect 240796 331294 240824 340068
rect 240888 340054 240994 340082
rect 241072 340054 241270 340082
rect 240784 331288 240836 331294
rect 240784 331230 240836 331236
rect 240888 331106 240916 340054
rect 241072 335646 241100 340054
rect 241060 335640 241112 335646
rect 241060 335582 241112 335588
rect 240612 331078 240916 331106
rect 240506 240136 240562 240145
rect 240506 240071 240562 240080
rect 240520 230518 240548 240071
rect 240508 230512 240560 230518
rect 240508 230454 240560 230460
rect 240506 220824 240562 220833
rect 240506 220759 240562 220768
rect 240520 211177 240548 220759
rect 240506 211168 240562 211177
rect 240506 211103 240562 211112
rect 240612 29102 240640 331078
rect 240692 331016 240744 331022
rect 240692 330958 240744 330964
rect 240704 299470 240732 330958
rect 240692 299464 240744 299470
rect 240692 299406 240744 299412
rect 240692 289876 240744 289882
rect 240692 289818 240744 289824
rect 240704 280158 240732 289818
rect 240692 280152 240744 280158
rect 240692 280094 240744 280100
rect 240692 270564 240744 270570
rect 240692 270506 240744 270512
rect 240704 240145 240732 270506
rect 240690 240136 240746 240145
rect 240690 240071 240746 240080
rect 240692 230512 240744 230518
rect 240692 230454 240744 230460
rect 240704 220833 240732 230454
rect 240690 220824 240746 220833
rect 240690 220759 240746 220768
rect 240690 211168 240746 211177
rect 240690 211103 240692 211112
rect 240744 211103 240746 211112
rect 240876 211132 240928 211138
rect 240692 211074 240744 211080
rect 240876 211074 240928 211080
rect 240888 201521 240916 211074
rect 240690 201512 240746 201521
rect 240690 201447 240746 201456
rect 240874 201512 240930 201521
rect 240874 201447 240930 201456
rect 240704 191826 240732 201447
rect 240692 191820 240744 191826
rect 240692 191762 240744 191768
rect 240876 191752 240928 191758
rect 240876 191694 240928 191700
rect 240888 182209 240916 191694
rect 240690 182200 240746 182209
rect 240690 182135 240746 182144
rect 240874 182200 240930 182209
rect 240874 182135 240930 182144
rect 240704 172514 240732 182135
rect 240692 172508 240744 172514
rect 240692 172450 240744 172456
rect 240876 172508 240928 172514
rect 240876 172450 240928 172456
rect 240888 162897 240916 172450
rect 240690 162888 240746 162897
rect 240690 162823 240746 162832
rect 240874 162888 240930 162897
rect 240874 162823 240930 162832
rect 240704 153202 240732 162823
rect 240692 153196 240744 153202
rect 240692 153138 240744 153144
rect 240876 153196 240928 153202
rect 240876 153138 240928 153144
rect 240888 143585 240916 153138
rect 240690 143576 240746 143585
rect 240690 143511 240692 143520
rect 240744 143511 240746 143520
rect 240874 143576 240930 143585
rect 240874 143511 240930 143520
rect 240692 143482 240744 143488
rect 240692 133952 240744 133958
rect 240692 133894 240744 133900
rect 240704 56574 240732 133894
rect 240692 56568 240744 56574
rect 240692 56510 240744 56516
rect 240692 47048 240744 47054
rect 240692 46990 240744 46996
rect 240704 46918 240732 46990
rect 240692 46912 240744 46918
rect 240692 46854 240744 46860
rect 240692 37392 240744 37398
rect 240692 37334 240744 37340
rect 240704 37262 240732 37334
rect 240692 37256 240744 37262
rect 240692 37198 240744 37204
rect 240600 29096 240652 29102
rect 240600 29038 240652 29044
rect 240600 28960 240652 28966
rect 240600 28902 240652 28908
rect 240416 6588 240468 6594
rect 240416 6530 240468 6536
rect 240324 6520 240376 6526
rect 240324 6462 240376 6468
rect 240138 5128 240194 5137
rect 240138 5063 240194 5072
rect 239404 4684 239456 4690
rect 239404 4626 239456 4632
rect 239588 4684 239640 4690
rect 239588 4626 239640 4632
rect 238852 4616 238904 4622
rect 238852 4558 238904 4564
rect 238864 4486 238892 4558
rect 238852 4480 238904 4486
rect 238852 4422 238904 4428
rect 239600 480 239628 4626
rect 240612 4622 240640 28902
rect 240692 18012 240744 18018
rect 240692 17954 240744 17960
rect 240704 7954 240732 17954
rect 241532 8022 241560 340068
rect 241716 338842 241744 340068
rect 241808 340054 242006 340082
rect 242176 340054 242282 340082
rect 242360 340054 242466 340082
rect 242544 340054 242742 340082
rect 241704 338836 241756 338842
rect 241704 338778 241756 338784
rect 241612 335640 241664 335646
rect 241612 335582 241664 335588
rect 241520 8016 241572 8022
rect 241520 7958 241572 7964
rect 240692 7948 240744 7954
rect 240692 7890 240744 7896
rect 241624 5438 241652 335582
rect 241808 6662 241836 340054
rect 242072 338836 242124 338842
rect 242072 338778 242124 338784
rect 241888 332036 241940 332042
rect 241888 331978 241940 331984
rect 241900 8090 241928 331978
rect 241888 8084 241940 8090
rect 241888 8026 241940 8032
rect 241796 6656 241848 6662
rect 241796 6598 241848 6604
rect 241612 5432 241664 5438
rect 241612 5374 241664 5380
rect 241980 5432 242032 5438
rect 241980 5374 242032 5380
rect 240600 4616 240652 4622
rect 240600 4558 240652 4564
rect 240784 4616 240836 4622
rect 240784 4558 240836 4564
rect 240796 480 240824 4558
rect 241992 480 242020 5374
rect 242084 5273 242112 338778
rect 242176 332042 242204 340054
rect 242360 335646 242388 340054
rect 242348 335640 242400 335646
rect 242348 335582 242400 335588
rect 242164 332036 242216 332042
rect 242164 331978 242216 331984
rect 242544 328574 242572 340054
rect 243004 338570 243032 340068
rect 243096 340054 243202 340082
rect 242992 338564 243044 338570
rect 242992 338506 243044 338512
rect 243096 335628 243124 340054
rect 243360 338972 243412 338978
rect 243360 338914 243412 338920
rect 243268 338564 243320 338570
rect 243268 338506 243320 338512
rect 242912 335600 243124 335628
rect 242532 328568 242584 328574
rect 242532 328510 242584 328516
rect 242256 328500 242308 328506
rect 242256 328442 242308 328448
rect 242268 19378 242296 328442
rect 242164 19372 242216 19378
rect 242164 19314 242216 19320
rect 242256 19372 242308 19378
rect 242256 19314 242308 19320
rect 242176 6730 242204 19314
rect 242164 6724 242216 6730
rect 242164 6666 242216 6672
rect 242912 5409 242940 335600
rect 243084 335504 243136 335510
rect 243084 335446 243136 335452
rect 243096 6866 243124 335446
rect 243280 8158 243308 338506
rect 243372 8226 243400 338914
rect 243360 8220 243412 8226
rect 243360 8162 243412 8168
rect 243268 8152 243320 8158
rect 243268 8094 243320 8100
rect 243084 6860 243136 6866
rect 243084 6802 243136 6808
rect 243464 6798 243492 340068
rect 243740 338978 243768 340068
rect 243832 340054 243938 340082
rect 244016 340054 244214 340082
rect 244384 340054 244490 340082
rect 244568 340054 244674 340082
rect 244752 340054 244950 340082
rect 243728 338972 243780 338978
rect 243728 338914 243780 338920
rect 243832 328506 243860 340054
rect 244016 335510 244044 340054
rect 244280 335640 244332 335646
rect 244280 335582 244332 335588
rect 244004 335504 244056 335510
rect 244004 335446 244056 335452
rect 243636 328500 243688 328506
rect 243636 328442 243688 328448
rect 243820 328500 243872 328506
rect 243820 328442 243872 328448
rect 243648 316690 243676 328442
rect 243556 316662 243676 316690
rect 243556 307034 243584 316662
rect 243556 307006 243676 307034
rect 243648 297378 243676 307006
rect 243556 297350 243676 297378
rect 243556 287722 243584 297350
rect 243556 287694 243676 287722
rect 243648 278066 243676 287694
rect 243556 278038 243676 278066
rect 243556 268410 243584 278038
rect 243556 268382 243676 268410
rect 243648 258754 243676 268382
rect 243556 258726 243676 258754
rect 243556 249098 243584 258726
rect 243556 249070 243676 249098
rect 243648 239442 243676 249070
rect 244186 240136 244242 240145
rect 244186 240071 244242 240080
rect 243556 239414 243676 239442
rect 243556 229786 243584 239414
rect 244200 234598 244228 240071
rect 244188 234592 244240 234598
rect 244188 234534 244240 234540
rect 243556 229758 243676 229786
rect 243648 220130 243676 229758
rect 243556 220102 243676 220130
rect 243556 210474 243584 220102
rect 243556 210446 243676 210474
rect 243648 200818 243676 210446
rect 243556 200790 243676 200818
rect 243556 191162 243584 200790
rect 244186 193216 244242 193225
rect 244186 193151 244242 193160
rect 243556 191134 243676 191162
rect 243648 181506 243676 191134
rect 244200 189514 244228 193151
rect 244188 189508 244240 189514
rect 244188 189450 244240 189456
rect 243556 181478 243676 181506
rect 243556 171850 243584 181478
rect 244186 173904 244242 173913
rect 244186 173839 244242 173848
rect 243556 171822 243676 171850
rect 243648 162194 243676 171822
rect 244200 164257 244228 173839
rect 244186 164248 244242 164257
rect 244186 164183 244188 164192
rect 244240 164183 244242 164192
rect 244188 164154 244240 164160
rect 243556 162166 243676 162194
rect 243556 152538 243584 162166
rect 244200 154601 244228 164154
rect 244186 154592 244242 154601
rect 244186 154527 244242 154536
rect 243556 152510 243676 152538
rect 243648 142882 243676 152510
rect 243556 142854 243676 142882
rect 243556 133226 243584 142854
rect 243556 133198 243676 133226
rect 243648 123570 243676 133198
rect 243556 123542 243676 123570
rect 243556 113914 243584 123542
rect 243556 113886 243676 113914
rect 243648 104258 243676 113886
rect 243556 104230 243676 104258
rect 243556 96778 243584 104230
rect 243556 96750 243676 96778
rect 243648 80170 243676 96750
rect 243636 80164 243688 80170
rect 243636 80106 243688 80112
rect 243544 80028 243596 80034
rect 243544 79970 243596 79976
rect 243556 77246 243584 79970
rect 243544 77240 243596 77246
rect 243544 77182 243596 77188
rect 243636 77240 243688 77246
rect 243636 77182 243688 77188
rect 243648 19378 243676 77182
rect 243544 19372 243596 19378
rect 243544 19314 243596 19320
rect 243636 19372 243688 19378
rect 243636 19314 243688 19320
rect 243452 6792 243504 6798
rect 243452 6734 243504 6740
rect 243556 5658 243584 19314
rect 243096 5630 243584 5658
rect 243096 5506 243124 5630
rect 243084 5500 243136 5506
rect 243084 5442 243136 5448
rect 243176 5500 243228 5506
rect 243176 5442 243228 5448
rect 242898 5400 242954 5409
rect 242898 5335 242954 5344
rect 242070 5264 242126 5273
rect 242070 5199 242126 5208
rect 243188 480 243216 5442
rect 244292 4758 244320 335582
rect 244384 334370 244412 340054
rect 244568 334490 244596 340054
rect 244556 334484 244608 334490
rect 244556 334426 244608 334432
rect 244384 334342 244596 334370
rect 244464 328500 244516 328506
rect 244464 328442 244516 328448
rect 244476 321638 244504 328442
rect 244464 321632 244516 321638
rect 244464 321574 244516 321580
rect 244464 321496 244516 321502
rect 244464 321438 244516 321444
rect 244476 318866 244504 321438
rect 244384 318838 244504 318866
rect 244384 317422 244412 318838
rect 244372 317416 244424 317422
rect 244372 317358 244424 317364
rect 244372 311500 244424 311506
rect 244372 311442 244424 311448
rect 244384 289882 244412 311442
rect 244372 289876 244424 289882
rect 244372 289818 244424 289824
rect 244464 289876 244516 289882
rect 244464 289818 244516 289824
rect 244476 278798 244504 289818
rect 244464 278792 244516 278798
rect 244464 278734 244516 278740
rect 244370 258088 244426 258097
rect 244370 258023 244372 258032
rect 244424 258023 244426 258032
rect 244372 257994 244424 258000
rect 244372 241596 244424 241602
rect 244372 241538 244424 241544
rect 244384 240145 244412 241538
rect 244370 240136 244426 240145
rect 244370 240071 244426 240080
rect 244372 234592 244424 234598
rect 244372 234534 244424 234540
rect 244384 217410 244412 234534
rect 244384 217382 244504 217410
rect 244476 202910 244504 217382
rect 244568 202978 244596 334342
rect 244648 278792 244700 278798
rect 244648 278734 244700 278740
rect 244660 258097 244688 278734
rect 244646 258088 244702 258097
rect 244646 258023 244702 258032
rect 244556 202972 244608 202978
rect 244556 202914 244608 202920
rect 244464 202904 244516 202910
rect 244464 202846 244516 202852
rect 244556 202836 244608 202842
rect 244556 202778 244608 202784
rect 244464 201544 244516 201550
rect 244464 201486 244516 201492
rect 244476 193225 244504 201486
rect 244462 193216 244518 193225
rect 244462 193151 244518 193160
rect 244464 173936 244516 173942
rect 244462 173904 244464 173913
rect 244516 173904 244518 173913
rect 244462 173839 244518 173848
rect 244370 164248 244426 164257
rect 244370 164183 244372 164192
rect 244424 164183 244426 164192
rect 244372 164154 244424 164160
rect 244462 154592 244518 154601
rect 244462 154527 244518 154536
rect 244476 147762 244504 154527
rect 244464 147756 244516 147762
rect 244464 147698 244516 147704
rect 244372 147620 244424 147626
rect 244372 147562 244424 147568
rect 244384 143546 244412 147562
rect 244372 143540 244424 143546
rect 244372 143482 244424 143488
rect 244464 143540 244516 143546
rect 244464 143482 244516 143488
rect 244476 138689 244504 143482
rect 244462 138680 244518 138689
rect 244462 138615 244518 138624
rect 244370 125624 244426 125633
rect 244370 125559 244426 125568
rect 244384 122806 244412 125559
rect 244372 122800 244424 122806
rect 244372 122742 244424 122748
rect 244464 113212 244516 113218
rect 244464 113154 244516 113160
rect 244476 113082 244504 113154
rect 244464 113076 244516 113082
rect 244464 113018 244516 113024
rect 244372 103624 244424 103630
rect 244372 103566 244424 103572
rect 244384 103494 244412 103566
rect 244372 103488 244424 103494
rect 244372 103430 244424 103436
rect 244464 85604 244516 85610
rect 244464 85546 244516 85552
rect 244476 84182 244504 85546
rect 244464 84176 244516 84182
rect 244464 84118 244516 84124
rect 244464 77240 244516 77246
rect 244464 77182 244516 77188
rect 244476 56574 244504 77182
rect 244464 56568 244516 56574
rect 244464 56510 244516 56516
rect 244372 46980 244424 46986
rect 244372 46922 244424 46928
rect 244384 41478 244412 46922
rect 244372 41472 244424 41478
rect 244372 41414 244424 41420
rect 244372 38616 244424 38622
rect 244372 38558 244424 38564
rect 244384 28914 244412 38558
rect 244384 28886 244504 28914
rect 244476 27606 244504 28886
rect 244464 27600 244516 27606
rect 244464 27542 244516 27548
rect 244464 18012 244516 18018
rect 244464 17954 244516 17960
rect 244476 12510 244504 17954
rect 244464 12504 244516 12510
rect 244464 12446 244516 12452
rect 244372 12436 244424 12442
rect 244372 12378 244424 12384
rect 244384 5370 244412 12378
rect 244568 8294 244596 202778
rect 244648 103488 244700 103494
rect 244648 103430 244700 103436
rect 244660 85610 244688 103430
rect 244648 85604 244700 85610
rect 244648 85546 244700 85552
rect 244556 8288 244608 8294
rect 244556 8230 244608 8236
rect 244752 6118 244780 340054
rect 245120 331242 245148 340068
rect 245212 340054 245410 340082
rect 245212 335646 245240 340054
rect 245200 335640 245252 335646
rect 245200 335582 245252 335588
rect 245120 331214 245240 331242
rect 245212 331106 245240 331214
rect 245028 331078 245240 331106
rect 245028 311930 245056 331078
rect 244936 311902 245056 311930
rect 244936 299538 244964 311902
rect 244924 299532 244976 299538
rect 244924 299474 244976 299480
rect 245016 299532 245068 299538
rect 245016 299474 245068 299480
rect 245028 298110 245056 299474
rect 245016 298104 245068 298110
rect 245016 298046 245068 298052
rect 244924 278792 244976 278798
rect 244924 278734 244976 278740
rect 244936 270502 244964 278734
rect 244924 270496 244976 270502
rect 244924 270438 244976 270444
rect 245108 270496 245160 270502
rect 245108 270438 245160 270444
rect 245120 259418 245148 270438
rect 244924 259412 244976 259418
rect 244924 259354 244976 259360
rect 245108 259412 245160 259418
rect 245108 259354 245160 259360
rect 244936 253042 244964 259354
rect 244936 253014 245056 253042
rect 245028 234666 245056 253014
rect 245016 234660 245068 234666
rect 245016 234602 245068 234608
rect 244924 234592 244976 234598
rect 244924 234534 244976 234540
rect 244936 227066 244964 234534
rect 244936 227038 245056 227066
rect 245028 212702 245056 227038
rect 245016 212696 245068 212702
rect 245016 212638 245068 212644
rect 245016 212492 245068 212498
rect 245016 212434 245068 212440
rect 245028 195294 245056 212434
rect 245016 195288 245068 195294
rect 245016 195230 245068 195236
rect 245016 183592 245068 183598
rect 245016 183534 245068 183540
rect 245028 178786 245056 183534
rect 245028 178758 245148 178786
rect 245120 173942 245148 178758
rect 244924 173936 244976 173942
rect 244924 173878 244976 173884
rect 245108 173936 245160 173942
rect 245108 173878 245160 173884
rect 244936 164393 244964 173878
rect 244922 164384 244978 164393
rect 244922 164319 244978 164328
rect 245014 164248 245070 164257
rect 245014 164183 245070 164192
rect 245028 157162 245056 164183
rect 244936 157134 245056 157162
rect 244936 147762 244964 157134
rect 244924 147756 244976 147762
rect 244924 147698 244976 147704
rect 244924 147620 244976 147626
rect 244924 147562 244976 147568
rect 244936 140758 244964 147562
rect 244924 140752 244976 140758
rect 244924 140694 244976 140700
rect 245108 131164 245160 131170
rect 245108 131106 245160 131112
rect 245120 121446 245148 131106
rect 245108 121440 245160 121446
rect 245108 121382 245160 121388
rect 245108 113144 245160 113150
rect 245108 113086 245160 113092
rect 245120 107030 245148 113086
rect 244924 107024 244976 107030
rect 244924 106966 244976 106972
rect 245108 107024 245160 107030
rect 245108 106966 245160 106972
rect 244936 99414 244964 106966
rect 244924 99408 244976 99414
rect 244924 99350 244976 99356
rect 245016 99340 245068 99346
rect 245016 99282 245068 99288
rect 245028 84182 245056 99282
rect 245016 84176 245068 84182
rect 245016 84118 245068 84124
rect 245108 84176 245160 84182
rect 245108 84118 245160 84124
rect 245120 75834 245148 84118
rect 245028 75806 245148 75834
rect 245028 58002 245056 75806
rect 244924 57996 244976 58002
rect 244924 57938 244976 57944
rect 245016 57996 245068 58002
rect 245016 57938 245068 57944
rect 244936 48346 244964 57938
rect 244924 48340 244976 48346
rect 244924 48282 244976 48288
rect 245016 48340 245068 48346
rect 245016 48282 245068 48288
rect 245028 28966 245056 48282
rect 244924 28960 244976 28966
rect 244924 28902 244976 28908
rect 245016 28960 245068 28966
rect 245016 28902 245068 28908
rect 244936 12510 244964 28902
rect 244924 12504 244976 12510
rect 244924 12446 244976 12452
rect 244832 12436 244884 12442
rect 244832 12378 244884 12384
rect 244844 7546 244872 12378
rect 244832 7540 244884 7546
rect 244832 7482 244884 7488
rect 244740 6112 244792 6118
rect 244740 6054 244792 6060
rect 245672 6050 245700 340068
rect 245752 335844 245804 335850
rect 245752 335786 245804 335792
rect 245660 6044 245712 6050
rect 245660 5986 245712 5992
rect 245764 5545 245792 335786
rect 245856 331294 245884 340068
rect 245948 340054 246146 340082
rect 246224 340054 246422 340082
rect 245948 335850 245976 340054
rect 245936 335844 245988 335850
rect 245936 335786 245988 335792
rect 246224 332194 246252 340054
rect 246132 332166 246252 332194
rect 245844 331288 245896 331294
rect 245844 331230 245896 331236
rect 246028 331152 246080 331158
rect 246028 331094 246080 331100
rect 245936 329180 245988 329186
rect 245936 329122 245988 329128
rect 245842 183560 245898 183569
rect 245842 183495 245898 183504
rect 245856 173942 245884 183495
rect 245844 173936 245896 173942
rect 245844 173878 245896 173884
rect 245844 133340 245896 133346
rect 245844 133282 245896 133288
rect 245856 124273 245884 133282
rect 245842 124264 245898 124273
rect 245842 124199 245898 124208
rect 245844 33856 245896 33862
rect 245844 33798 245896 33804
rect 245856 19378 245884 33798
rect 245844 19372 245896 19378
rect 245844 19314 245896 19320
rect 245948 5982 245976 329122
rect 246040 280158 246068 331094
rect 246132 329186 246160 332166
rect 246212 332104 246264 332110
rect 246212 332046 246264 332052
rect 246120 329180 246172 329186
rect 246120 329122 246172 329128
rect 246028 280152 246080 280158
rect 246028 280094 246080 280100
rect 246028 270564 246080 270570
rect 246028 270506 246080 270512
rect 246040 183569 246068 270506
rect 246026 183560 246082 183569
rect 246026 183495 246082 183504
rect 246028 173936 246080 173942
rect 246028 173878 246080 173884
rect 246040 143546 246068 173878
rect 246028 143540 246080 143546
rect 246028 143482 246080 143488
rect 246026 124264 246082 124273
rect 246026 124199 246082 124208
rect 246040 87038 246068 124199
rect 246028 87032 246080 87038
rect 246028 86974 246080 86980
rect 246120 86896 246172 86902
rect 246120 86838 246172 86844
rect 246132 77382 246160 86838
rect 246120 77376 246172 77382
rect 246120 77318 246172 77324
rect 246028 74588 246080 74594
rect 246028 74530 246080 74536
rect 246040 33862 246068 74530
rect 246028 33856 246080 33862
rect 246028 33798 246080 33804
rect 246028 19372 246080 19378
rect 246028 19314 246080 19320
rect 246040 7478 246068 19314
rect 246028 7472 246080 7478
rect 246028 7414 246080 7420
rect 245936 5976 245988 5982
rect 245936 5918 245988 5924
rect 245750 5536 245806 5545
rect 245750 5471 245806 5480
rect 244372 5364 244424 5370
rect 244372 5306 244424 5312
rect 244648 5364 244700 5370
rect 244648 5306 244700 5312
rect 244280 4752 244332 4758
rect 244280 4694 244332 4700
rect 244660 2802 244688 5306
rect 245568 4752 245620 4758
rect 245568 4694 245620 4700
rect 244476 2774 244688 2802
rect 244476 2666 244504 2774
rect 244384 2638 244504 2666
rect 244384 480 244412 2638
rect 245580 480 245608 4694
rect 246224 4486 246252 332046
rect 246592 331276 246620 340068
rect 246684 340054 246882 340082
rect 247158 340054 247264 340082
rect 247342 340054 247448 340082
rect 246684 332110 246712 340054
rect 247040 335708 247092 335714
rect 247040 335650 247092 335656
rect 246672 332104 246724 332110
rect 246672 332046 246724 332052
rect 246592 331248 246712 331276
rect 246684 331106 246712 331248
rect 246500 331078 246712 331106
rect 246500 311930 246528 331078
rect 246408 311902 246528 311930
rect 246408 309126 246436 311902
rect 246396 309120 246448 309126
rect 246396 309062 246448 309068
rect 246488 309052 246540 309058
rect 246488 308994 246540 309000
rect 246500 299470 246528 308994
rect 246396 299464 246448 299470
rect 246396 299406 246448 299412
rect 246488 299464 246540 299470
rect 246488 299406 246540 299412
rect 246408 288386 246436 299406
rect 246396 288380 246448 288386
rect 246396 288322 246448 288328
rect 246488 278792 246540 278798
rect 246488 278734 246540 278740
rect 246500 272610 246528 278734
rect 246488 272604 246540 272610
rect 246488 272546 246540 272552
rect 246764 272604 246816 272610
rect 246764 272546 246816 272552
rect 246776 267889 246804 272546
rect 246486 267880 246542 267889
rect 246486 267815 246542 267824
rect 246762 267880 246818 267889
rect 246762 267815 246818 267824
rect 246500 267753 246528 267815
rect 246302 267744 246358 267753
rect 246302 267679 246358 267688
rect 246486 267744 246542 267753
rect 246486 267679 246542 267688
rect 246316 258126 246344 267679
rect 246304 258120 246356 258126
rect 246304 258062 246356 258068
rect 246396 258120 246448 258126
rect 246396 258062 246448 258068
rect 246408 253178 246436 258062
rect 246316 253150 246436 253178
rect 246316 248402 246344 253150
rect 246304 248396 246356 248402
rect 246304 248338 246356 248344
rect 246396 238808 246448 238814
rect 246396 238750 246448 238756
rect 246408 234666 246436 238750
rect 246396 234660 246448 234666
rect 246396 234602 246448 234608
rect 246488 234524 246540 234530
rect 246488 234466 246540 234472
rect 246500 217462 246528 234466
rect 246488 217456 246540 217462
rect 246488 217398 246540 217404
rect 246396 209840 246448 209846
rect 246396 209782 246448 209788
rect 246408 205698 246436 209782
rect 246396 205692 246448 205698
rect 246396 205634 246448 205640
rect 246488 205556 246540 205562
rect 246488 205498 246540 205504
rect 246500 198098 246528 205498
rect 246500 198070 246620 198098
rect 246592 193254 246620 198070
rect 246396 193248 246448 193254
rect 246394 193216 246396 193225
rect 246580 193248 246632 193254
rect 246448 193216 246450 193225
rect 246394 193151 246450 193160
rect 246578 193216 246580 193225
rect 246632 193216 246634 193225
rect 246578 193151 246634 193160
rect 246592 186266 246620 193151
rect 246500 186238 246620 186266
rect 246500 178786 246528 186238
rect 246500 178758 246620 178786
rect 246592 173942 246620 178758
rect 246396 173936 246448 173942
rect 246396 173878 246448 173884
rect 246580 173936 246632 173942
rect 246580 173878 246632 173884
rect 246408 169402 246436 173878
rect 246408 169374 246528 169402
rect 246500 154737 246528 169374
rect 246486 154728 246542 154737
rect 246486 154663 246542 154672
rect 246394 154592 246450 154601
rect 246394 154527 246450 154536
rect 246408 143614 246436 154527
rect 246396 143608 246448 143614
rect 246396 143550 246448 143556
rect 246396 142180 246448 142186
rect 246396 142122 246448 142128
rect 246408 142050 246436 142122
rect 246396 142044 246448 142050
rect 246396 141986 246448 141992
rect 246396 124228 246448 124234
rect 246396 124170 246448 124176
rect 246408 114458 246436 124170
rect 246408 114430 246620 114458
rect 246592 104922 246620 114430
rect 246488 104916 246540 104922
rect 246488 104858 246540 104864
rect 246580 104916 246632 104922
rect 246580 104858 246632 104864
rect 246500 99482 246528 104858
rect 246488 99476 246540 99482
rect 246488 99418 246540 99424
rect 246304 95192 246356 95198
rect 246304 95134 246356 95140
rect 246316 85610 246344 95134
rect 246304 85604 246356 85610
rect 246304 85546 246356 85552
rect 246396 85604 246448 85610
rect 246396 85546 246448 85552
rect 246408 77625 246436 85546
rect 246394 77616 246450 77625
rect 246394 77551 246450 77560
rect 246394 77344 246450 77353
rect 246394 77279 246450 77288
rect 246408 71074 246436 77279
rect 246408 71046 246620 71074
rect 246592 57934 246620 71046
rect 246580 57928 246632 57934
rect 246580 57870 246632 57876
rect 246488 48340 246540 48346
rect 246488 48282 246540 48288
rect 246500 18018 246528 48282
rect 246946 40488 247002 40497
rect 246946 40423 247002 40432
rect 246960 40361 246988 40423
rect 246946 40352 247002 40361
rect 246946 40287 247002 40296
rect 246304 18012 246356 18018
rect 246304 17954 246356 17960
rect 246488 18012 246540 18018
rect 246488 17954 246540 17960
rect 246316 8208 246344 17954
rect 246316 8180 246436 8208
rect 246408 7410 246436 8180
rect 246396 7404 246448 7410
rect 246396 7346 246448 7352
rect 246764 4616 246816 4622
rect 246764 4558 246816 4564
rect 246212 4480 246264 4486
rect 246212 4422 246264 4428
rect 246776 480 246804 4558
rect 247052 4418 247080 335650
rect 247236 5914 247264 340054
rect 247420 7342 247448 340054
rect 247500 335640 247552 335646
rect 247500 335582 247552 335588
rect 247408 7336 247460 7342
rect 247408 7278 247460 7284
rect 247512 7274 247540 335582
rect 247500 7268 247552 7274
rect 247500 7210 247552 7216
rect 247224 5908 247276 5914
rect 247224 5850 247276 5856
rect 247604 4554 247632 340068
rect 247696 340054 247894 340082
rect 247972 340054 248078 340082
rect 248156 340054 248354 340082
rect 247696 5846 247724 340054
rect 247972 335646 248000 340054
rect 248156 335714 248184 340054
rect 248144 335708 248196 335714
rect 248144 335650 248196 335656
rect 248420 335708 248472 335714
rect 248420 335650 248472 335656
rect 247960 335640 248012 335646
rect 247960 335582 248012 335588
rect 247684 5840 247736 5846
rect 247684 5782 247736 5788
rect 247592 4548 247644 4554
rect 247592 4490 247644 4496
rect 247960 4548 248012 4554
rect 247960 4490 248012 4496
rect 247040 4412 247092 4418
rect 247040 4354 247092 4360
rect 247972 480 248000 4490
rect 248432 4282 248460 335650
rect 248512 335572 248564 335578
rect 248512 335514 248564 335520
rect 248524 5710 248552 335514
rect 248616 5778 248644 340068
rect 248696 335640 248748 335646
rect 248696 335582 248748 335588
rect 248708 7138 248736 335582
rect 248800 7206 248828 340068
rect 248892 340054 249090 340082
rect 249168 340054 249366 340082
rect 249444 340054 249550 340082
rect 248892 335714 248920 340054
rect 248880 335708 248932 335714
rect 248880 335650 248932 335656
rect 249168 335578 249196 340054
rect 249444 335646 249472 340054
rect 249432 335640 249484 335646
rect 249432 335582 249484 335588
rect 249156 335572 249208 335578
rect 249156 335514 249208 335520
rect 249706 87000 249762 87009
rect 249706 86935 249708 86944
rect 249760 86935 249762 86944
rect 249708 86906 249760 86912
rect 248788 7200 248840 7206
rect 248788 7142 248840 7148
rect 248696 7132 248748 7138
rect 248696 7074 248748 7080
rect 248604 5772 248656 5778
rect 248604 5714 248656 5720
rect 248512 5704 248564 5710
rect 248512 5646 248564 5652
rect 249812 4282 249840 340068
rect 249892 335708 249944 335714
rect 249892 335650 249944 335656
rect 249904 4350 249932 335650
rect 249984 335572 250036 335578
rect 249984 335514 250036 335520
rect 249996 5574 250024 335514
rect 250088 5642 250116 340068
rect 250168 335640 250220 335646
rect 250168 335582 250220 335588
rect 250180 7002 250208 335582
rect 250272 7070 250300 340068
rect 250364 340054 250562 340082
rect 250640 340054 250838 340082
rect 250916 340054 251022 340082
rect 251192 340054 251298 340082
rect 250364 335714 250392 340054
rect 250352 335708 250404 335714
rect 250352 335650 250404 335656
rect 250640 335578 250668 340054
rect 250916 335646 250944 340054
rect 250904 335640 250956 335646
rect 250904 335582 250956 335588
rect 250628 335572 250680 335578
rect 250628 335514 250680 335520
rect 250260 7064 250312 7070
rect 250260 7006 250312 7012
rect 250168 6996 250220 7002
rect 250168 6938 250220 6944
rect 250076 5636 250128 5642
rect 250076 5578 250128 5584
rect 249984 5568 250036 5574
rect 249984 5510 250036 5516
rect 251192 4826 251220 340054
rect 251364 335708 251416 335714
rect 251364 335650 251416 335656
rect 251376 5030 251404 335650
rect 251456 335572 251508 335578
rect 251456 335514 251508 335520
rect 251468 5302 251496 335514
rect 251456 5296 251508 5302
rect 251456 5238 251508 5244
rect 251364 5024 251416 5030
rect 251364 4966 251416 4972
rect 251560 4894 251588 340068
rect 251640 335640 251692 335646
rect 251640 335582 251692 335588
rect 251652 5098 251680 335582
rect 251640 5092 251692 5098
rect 251640 5034 251692 5040
rect 251744 4962 251772 340068
rect 251836 340054 252034 340082
rect 252112 340054 252310 340082
rect 252388 340054 252494 340082
rect 251836 335714 251864 340054
rect 251824 335708 251876 335714
rect 251824 335650 251876 335656
rect 252112 335646 252140 340054
rect 252100 335640 252152 335646
rect 252100 335582 252152 335588
rect 252388 335578 252416 340054
rect 252652 335708 252704 335714
rect 252652 335650 252704 335656
rect 252560 335640 252612 335646
rect 252560 335582 252612 335588
rect 252376 335572 252428 335578
rect 252376 335514 252428 335520
rect 252100 86964 252152 86970
rect 252100 86906 252152 86912
rect 252112 86873 252140 86906
rect 252098 86864 252154 86873
rect 252098 86799 252154 86808
rect 251732 4956 251784 4962
rect 251732 4898 251784 4904
rect 251548 4888 251600 4894
rect 251548 4830 251600 4836
rect 251180 4820 251232 4826
rect 251180 4762 251232 4768
rect 252572 4690 252600 335582
rect 252664 5574 252692 335650
rect 252652 5568 252704 5574
rect 252652 5510 252704 5516
rect 252756 5166 252784 340068
rect 252848 340054 253046 340082
rect 253124 340054 253230 340082
rect 253308 340054 253506 340082
rect 253676 340054 253782 340082
rect 253966 340054 254072 340082
rect 252848 5234 252876 340054
rect 253124 335646 253152 340054
rect 253308 335714 253336 340054
rect 253296 335708 253348 335714
rect 253296 335650 253348 335656
rect 253112 335640 253164 335646
rect 253112 335582 253164 335588
rect 253676 328506 253704 340054
rect 253112 328500 253164 328506
rect 253112 328442 253164 328448
rect 253664 328500 253716 328506
rect 253664 328442 253716 328448
rect 253124 311930 253152 328442
rect 253032 311902 253152 311930
rect 253032 311794 253060 311902
rect 253032 311766 253152 311794
rect 253124 309126 253152 311766
rect 253112 309120 253164 309126
rect 253112 309062 253164 309068
rect 253204 309120 253256 309126
rect 253204 309062 253256 309068
rect 253216 289882 253244 309062
rect 253020 289876 253072 289882
rect 253020 289818 253072 289824
rect 253204 289876 253256 289882
rect 253204 289818 253256 289824
rect 253032 269113 253060 289818
rect 253018 269104 253074 269113
rect 253018 269039 253074 269048
rect 253110 268968 253166 268977
rect 253110 268903 253166 268912
rect 253124 254046 253152 268903
rect 253112 254040 253164 254046
rect 253112 253982 253164 253988
rect 253020 253904 253072 253910
rect 253020 253846 253072 253852
rect 253032 241534 253060 253846
rect 253020 241528 253072 241534
rect 253020 241470 253072 241476
rect 253112 241528 253164 241534
rect 253112 241470 253164 241476
rect 253124 230586 253152 241470
rect 253020 230580 253072 230586
rect 253020 230522 253072 230528
rect 253112 230580 253164 230586
rect 253112 230522 253164 230528
rect 253032 230489 253060 230522
rect 253018 230480 253074 230489
rect 253018 230415 253074 230424
rect 253294 230480 253350 230489
rect 253294 230415 253350 230424
rect 253308 220862 253336 230415
rect 253112 220856 253164 220862
rect 253112 220798 253164 220804
rect 253296 220856 253348 220862
rect 253296 220798 253348 220804
rect 253124 217546 253152 220798
rect 253124 217518 253244 217546
rect 253216 211177 253244 217518
rect 253018 211168 253074 211177
rect 253018 211103 253074 211112
rect 253202 211168 253258 211177
rect 253202 211103 253258 211112
rect 253032 202910 253060 211103
rect 253020 202904 253072 202910
rect 253020 202846 253072 202852
rect 253112 202904 253164 202910
rect 253112 202846 253164 202852
rect 253124 191894 253152 202846
rect 253020 191888 253072 191894
rect 253020 191830 253072 191836
rect 253112 191888 253164 191894
rect 253112 191830 253164 191836
rect 253032 186946 253060 191830
rect 253032 186918 253152 186946
rect 253124 177426 253152 186918
rect 253032 177398 253152 177426
rect 253032 172582 253060 177398
rect 252928 172576 252980 172582
rect 252928 172518 252980 172524
rect 253020 172576 253072 172582
rect 253020 172518 253072 172524
rect 252940 164286 252968 172518
rect 252928 164280 252980 164286
rect 252928 164222 252980 164228
rect 253020 164280 253072 164286
rect 253020 164222 253072 164228
rect 253032 161430 253060 164222
rect 253020 161424 253072 161430
rect 253020 161366 253072 161372
rect 253020 151836 253072 151842
rect 253020 151778 253072 151784
rect 253032 151706 253060 151778
rect 253020 151700 253072 151706
rect 253020 151642 253072 151648
rect 253204 142248 253256 142254
rect 253204 142190 253256 142196
rect 253216 140758 253244 142190
rect 253204 140752 253256 140758
rect 253204 140694 253256 140700
rect 253204 131164 253256 131170
rect 253204 131106 253256 131112
rect 253216 122890 253244 131106
rect 253032 122862 253244 122890
rect 253032 122806 253060 122862
rect 253020 122800 253072 122806
rect 253020 122742 253072 122748
rect 253204 108384 253256 108390
rect 253204 108326 253256 108332
rect 253216 103494 253244 108326
rect 253204 103488 253256 103494
rect 253204 103430 253256 103436
rect 253204 95192 253256 95198
rect 253204 95134 253256 95140
rect 253216 85678 253244 95134
rect 253204 85672 253256 85678
rect 253204 85614 253256 85620
rect 253020 84244 253072 84250
rect 253020 84186 253072 84192
rect 253032 84114 253060 84186
rect 253020 84108 253072 84114
rect 253020 84050 253072 84056
rect 253112 84108 253164 84114
rect 253112 84050 253164 84056
rect 253124 74594 253152 84050
rect 253112 74588 253164 74594
rect 253112 74530 253164 74536
rect 253296 74452 253348 74458
rect 253296 74394 253348 74400
rect 253308 73166 253336 74394
rect 253296 73160 253348 73166
rect 253296 73102 253348 73108
rect 253204 63572 253256 63578
rect 253204 63514 253256 63520
rect 253216 63458 253244 63514
rect 253216 63430 253336 63458
rect 253308 63322 253336 63430
rect 253308 63294 253428 63322
rect 253400 55162 253428 63294
rect 253308 55134 253428 55162
rect 253308 50386 253336 55134
rect 253020 50380 253072 50386
rect 253020 50322 253072 50328
rect 253296 50380 253348 50386
rect 253296 50322 253348 50328
rect 253032 45558 253060 50322
rect 253020 45552 253072 45558
rect 253020 45494 253072 45500
rect 252928 40724 252980 40730
rect 252928 40666 252980 40672
rect 252940 35902 252968 40666
rect 252928 35896 252980 35902
rect 252928 35838 252980 35844
rect 253020 26308 253072 26314
rect 253020 26250 253072 26256
rect 253032 26194 253060 26250
rect 253110 26208 253166 26217
rect 253032 26166 253110 26194
rect 253110 26143 253166 26152
rect 253294 26208 253350 26217
rect 253294 26143 253350 26152
rect 253308 17882 253336 26143
rect 253112 17876 253164 17882
rect 253112 17818 253164 17824
rect 253296 17876 253348 17882
rect 253296 17818 253348 17824
rect 253124 8378 253152 17818
rect 252940 8350 253152 8378
rect 252940 8294 252968 8350
rect 252928 8288 252980 8294
rect 252928 8230 252980 8236
rect 254044 5506 254072 340054
rect 254308 335708 254360 335714
rect 254308 335650 254360 335656
rect 254124 335640 254176 335646
rect 254124 335582 254176 335588
rect 254032 5500 254084 5506
rect 254032 5442 254084 5448
rect 252836 5228 252888 5234
rect 252836 5170 252888 5176
rect 252744 5160 252796 5166
rect 252744 5102 252796 5108
rect 252560 4684 252612 4690
rect 252560 4626 252612 4632
rect 254136 4554 254164 335582
rect 254320 4758 254348 335650
rect 254412 5370 254440 340190
rect 254504 335714 254532 340068
rect 254596 340054 254702 340082
rect 254780 340054 254978 340082
rect 255056 340054 255254 340082
rect 255332 340054 255438 340082
rect 255608 340054 255714 340082
rect 255884 340054 255990 340082
rect 256068 340054 256174 340082
rect 256252 340054 256450 340082
rect 254492 335708 254544 335714
rect 254492 335650 254544 335656
rect 254490 29472 254546 29481
rect 254490 29407 254546 29416
rect 254504 29073 254532 29407
rect 254490 29064 254546 29073
rect 254490 28999 254546 29008
rect 254400 5364 254452 5370
rect 254400 5306 254452 5312
rect 254308 4752 254360 4758
rect 254308 4694 254360 4700
rect 254596 4622 254624 340054
rect 254780 335646 254808 340054
rect 254768 335640 254820 335646
rect 254768 335582 254820 335588
rect 255056 328681 255084 340054
rect 255042 328672 255098 328681
rect 255042 328607 255098 328616
rect 254674 328536 254730 328545
rect 254674 328471 254730 328480
rect 254688 328438 254716 328471
rect 254676 328432 254728 328438
rect 254676 328374 254728 328380
rect 254860 318844 254912 318850
rect 254860 318786 254912 318792
rect 254872 309126 254900 318786
rect 254676 309120 254728 309126
rect 254676 309062 254728 309068
rect 254860 309120 254912 309126
rect 254860 309062 254912 309068
rect 254688 299538 254716 309062
rect 254676 299532 254728 299538
rect 254676 299474 254728 299480
rect 254860 299396 254912 299402
rect 254860 299338 254912 299344
rect 254872 298058 254900 299338
rect 254872 298030 254992 298058
rect 254964 288454 254992 298030
rect 254860 288448 254912 288454
rect 254860 288390 254912 288396
rect 254952 288448 255004 288454
rect 254952 288390 255004 288396
rect 254872 280226 254900 288390
rect 254768 280220 254820 280226
rect 254768 280162 254820 280168
rect 254860 280220 254912 280226
rect 254860 280162 254912 280168
rect 254780 263650 254808 280162
rect 254688 263622 254808 263650
rect 254688 263514 254716 263622
rect 254688 263486 254808 263514
rect 254780 244338 254808 263486
rect 254688 244310 254808 244338
rect 254688 244202 254716 244310
rect 254688 244174 254808 244202
rect 254780 225026 254808 244174
rect 254688 224998 254808 225026
rect 254688 224890 254716 224998
rect 254688 224862 254808 224890
rect 254780 205714 254808 224862
rect 254688 205686 254808 205714
rect 254688 205578 254716 205686
rect 254688 205550 254808 205578
rect 254780 186402 254808 205550
rect 254688 186374 254808 186402
rect 254688 186266 254716 186374
rect 254688 186238 254808 186266
rect 254780 164393 254808 186238
rect 254766 164384 254822 164393
rect 254766 164319 254822 164328
rect 254766 164248 254822 164257
rect 254766 164183 254822 164192
rect 254780 143562 254808 164183
rect 254688 143546 254808 143562
rect 254676 143540 254808 143546
rect 254728 143534 254808 143540
rect 254860 143540 254912 143546
rect 254676 143482 254728 143488
rect 254860 143482 254912 143488
rect 254872 133906 254900 143482
rect 254872 133878 254992 133906
rect 254964 127650 254992 133878
rect 254780 127622 254992 127650
rect 254780 122806 254808 127622
rect 254768 122800 254820 122806
rect 254768 122742 254820 122748
rect 254676 104916 254728 104922
rect 254676 104858 254728 104864
rect 254688 95266 254716 104858
rect 254676 95260 254728 95266
rect 254676 95202 254728 95208
rect 254768 95260 254820 95266
rect 254768 95202 254820 95208
rect 254780 75886 254808 95202
rect 254768 75880 254820 75886
rect 254768 75822 254820 75828
rect 254952 69692 255004 69698
rect 254952 69634 255004 69640
rect 254964 64954 254992 69634
rect 254872 64926 254992 64954
rect 254872 63510 254900 64926
rect 254860 63504 254912 63510
rect 254860 63446 254912 63452
rect 254768 53848 254820 53854
rect 254768 53790 254820 53796
rect 254780 45558 254808 53790
rect 254768 45552 254820 45558
rect 254768 45494 254820 45500
rect 254768 45416 254820 45422
rect 254768 45358 254820 45364
rect 254780 29050 254808 45358
rect 254780 29022 254900 29050
rect 254872 28948 254900 29022
rect 254780 28920 254900 28948
rect 254584 4616 254636 4622
rect 254584 4558 254636 4564
rect 254124 4548 254176 4554
rect 254124 4490 254176 4496
rect 250352 4480 250404 4486
rect 250352 4422 250404 4428
rect 249892 4344 249944 4350
rect 249892 4286 249944 4292
rect 248420 4276 248472 4282
rect 248420 4218 248472 4224
rect 249800 4276 249852 4282
rect 249800 4218 249852 4224
rect 249156 4208 249208 4214
rect 249156 4150 249208 4156
rect 249168 480 249196 4150
rect 250364 480 250392 4422
rect 251456 4412 251508 4418
rect 251456 4354 251508 4360
rect 251468 480 251496 4354
rect 252652 4344 252704 4350
rect 252652 4286 252704 4292
rect 252664 480 252692 4286
rect 253848 4276 253900 4282
rect 253848 4218 253900 4224
rect 253860 480 253888 4218
rect 254780 4214 254808 28920
rect 255044 5500 255096 5506
rect 255044 5442 255096 5448
rect 254768 4208 254820 4214
rect 254768 4150 254820 4156
rect 255056 480 255084 5442
rect 255332 4486 255360 340054
rect 255504 335708 255556 335714
rect 255504 335650 255556 335656
rect 255320 4480 255372 4486
rect 255320 4422 255372 4428
rect 255516 4282 255544 335650
rect 255608 4418 255636 340054
rect 255780 335640 255832 335646
rect 255780 335582 255832 335588
rect 255792 5506 255820 335582
rect 255780 5500 255832 5506
rect 255780 5442 255832 5448
rect 255596 4412 255648 4418
rect 255596 4354 255648 4360
rect 255884 4350 255912 340054
rect 256068 335714 256096 340054
rect 256056 335708 256108 335714
rect 256056 335650 256108 335656
rect 256252 335646 256280 340054
rect 256240 335640 256292 335646
rect 256240 335582 256292 335588
rect 256712 334150 256740 340068
rect 256700 334144 256752 334150
rect 256700 334086 256752 334092
rect 256896 333418 256924 340068
rect 256712 333390 256924 333418
rect 256988 340054 257186 340082
rect 257264 340054 257462 340082
rect 257540 340054 257646 340082
rect 257724 340054 257922 340082
rect 256712 328545 256740 333390
rect 256988 333282 257016 340054
rect 257264 335560 257292 340054
rect 257344 335640 257396 335646
rect 257344 335582 257396 335588
rect 256804 333254 257016 333282
rect 257172 335532 257292 335560
rect 256698 328536 256754 328545
rect 256698 328471 256754 328480
rect 256804 326194 256832 333254
rect 257172 333146 257200 335532
rect 257252 334144 257304 334150
rect 257252 334086 257304 334092
rect 256988 333118 257200 333146
rect 256988 326262 257016 333118
rect 257066 328536 257122 328545
rect 257066 328471 257122 328480
rect 257080 327078 257108 328471
rect 257068 327072 257120 327078
rect 257068 327014 257120 327020
rect 256976 326256 257028 326262
rect 256976 326198 257028 326204
rect 256792 326188 256844 326194
rect 256792 326130 256844 326136
rect 257160 317484 257212 317490
rect 257160 317426 257212 317432
rect 257172 309126 257200 317426
rect 257068 309120 257120 309126
rect 257068 309062 257120 309068
rect 257160 309120 257212 309126
rect 257160 309062 257212 309068
rect 257080 302938 257108 309062
rect 257068 302932 257120 302938
rect 257068 302874 257120 302880
rect 257160 294500 257212 294506
rect 257160 294442 257212 294448
rect 257172 280158 257200 294442
rect 257160 280152 257212 280158
rect 257160 280094 257212 280100
rect 257160 278792 257212 278798
rect 257160 278734 257212 278740
rect 257080 259486 257108 259517
rect 257172 259486 257200 278734
rect 257068 259480 257120 259486
rect 256988 259428 257068 259434
rect 256988 259422 257120 259428
rect 257160 259480 257212 259486
rect 257160 259422 257212 259428
rect 256988 259406 257108 259422
rect 256988 251258 257016 259406
rect 256976 251252 257028 251258
rect 256976 251194 257028 251200
rect 256976 249824 257028 249830
rect 256976 249766 257028 249772
rect 256988 243930 257016 249766
rect 256988 243902 257108 243930
rect 257080 230518 257108 243902
rect 257068 230512 257120 230518
rect 257160 230512 257212 230518
rect 257120 230460 257160 230466
rect 257068 230454 257212 230460
rect 257080 230438 257200 230454
rect 257080 225010 257108 230438
rect 257068 225004 257120 225010
rect 257068 224946 257120 224952
rect 257160 224936 257212 224942
rect 257160 224878 257212 224884
rect 257172 202978 257200 224878
rect 257160 202972 257212 202978
rect 257160 202914 257212 202920
rect 257068 202904 257120 202910
rect 257068 202846 257120 202852
rect 257080 191842 257108 202846
rect 257080 191814 257200 191842
rect 257172 186454 257200 191814
rect 257160 186448 257212 186454
rect 257160 186390 257212 186396
rect 257068 186312 257120 186318
rect 257068 186254 257120 186260
rect 257080 172582 257108 186254
rect 256976 172576 257028 172582
rect 256976 172518 257028 172524
rect 257068 172576 257120 172582
rect 257068 172518 257120 172524
rect 256988 164286 257016 172518
rect 256976 164280 257028 164286
rect 256976 164222 257028 164228
rect 257068 164280 257120 164286
rect 257068 164222 257120 164228
rect 257080 161430 257108 164222
rect 257068 161424 257120 161430
rect 257068 161366 257120 161372
rect 257264 153270 257292 334086
rect 257356 326380 257384 335582
rect 257540 326482 257568 340054
rect 257724 335646 257752 340054
rect 257712 335640 257764 335646
rect 257712 335582 257764 335588
rect 258184 335510 258212 340068
rect 258276 340054 258382 340082
rect 258172 335504 258224 335510
rect 258172 335446 258224 335452
rect 258276 330750 258304 340054
rect 258644 335646 258672 340068
rect 258934 340054 259040 340082
rect 258724 338904 258776 338910
rect 258724 338846 258776 338852
rect 258632 335640 258684 335646
rect 258632 335582 258684 335588
rect 258632 335436 258684 335442
rect 258632 335378 258684 335384
rect 258264 330744 258316 330750
rect 258264 330686 258316 330692
rect 258644 328438 258672 335378
rect 258632 328432 258684 328438
rect 258632 328374 258684 328380
rect 257540 326454 258028 326482
rect 257356 326352 257936 326380
rect 257712 326256 257764 326262
rect 257712 326198 257764 326204
rect 257252 153264 257304 153270
rect 257252 153206 257304 153212
rect 257252 153128 257304 153134
rect 257252 153070 257304 153076
rect 256976 142180 257028 142186
rect 256976 142122 257028 142128
rect 256988 124273 257016 142122
rect 256974 124264 257030 124273
rect 256974 124199 257030 124208
rect 257158 124264 257214 124273
rect 257158 124199 257214 124208
rect 257172 122806 257200 124199
rect 257160 122800 257212 122806
rect 257160 122742 257212 122748
rect 257160 113212 257212 113218
rect 257160 113154 257212 113160
rect 257172 109698 257200 113154
rect 257080 109670 257200 109698
rect 257080 100042 257108 109670
rect 257080 100014 257200 100042
rect 257172 95198 257200 100014
rect 257160 95192 257212 95198
rect 257160 95134 257212 95140
rect 257068 85604 257120 85610
rect 257068 85546 257120 85552
rect 257080 74594 257108 85546
rect 257068 74588 257120 74594
rect 257068 74530 257120 74536
rect 257160 74588 257212 74594
rect 257160 74530 257212 74536
rect 257172 47122 257200 74530
rect 257160 47116 257212 47122
rect 257160 47058 257212 47064
rect 257160 46980 257212 46986
rect 257160 46922 257212 46928
rect 257172 45558 257200 46922
rect 257160 45552 257212 45558
rect 257160 45494 257212 45500
rect 256606 40624 256662 40633
rect 256606 40559 256662 40568
rect 256620 40225 256648 40559
rect 256606 40216 256662 40225
rect 256606 40151 256662 40160
rect 257160 27668 257212 27674
rect 257160 27610 257212 27616
rect 256240 5500 256292 5506
rect 256240 5442 256292 5448
rect 255872 4344 255924 4350
rect 255872 4286 255924 4292
rect 255504 4276 255556 4282
rect 255504 4218 255556 4224
rect 256252 480 256280 5442
rect 257172 5386 257200 27610
rect 257264 5506 257292 153070
rect 257344 151836 257396 151842
rect 257344 151778 257396 151784
rect 257356 142186 257384 151778
rect 257344 142180 257396 142186
rect 257344 142122 257396 142128
rect 257252 5500 257304 5506
rect 257252 5442 257304 5448
rect 257724 5438 257752 326198
rect 257804 326188 257856 326194
rect 257804 326130 257856 326136
rect 257816 5506 257844 326130
rect 257804 5500 257856 5506
rect 257804 5442 257856 5448
rect 257712 5432 257764 5438
rect 257172 5358 257476 5386
rect 257712 5374 257764 5380
rect 257448 480 257476 5358
rect 257908 5302 257936 326352
rect 258000 5370 258028 326454
rect 258736 326398 258764 338846
rect 259012 335594 259040 340054
rect 259104 338910 259132 340068
rect 259288 340054 259394 340082
rect 259670 340054 259776 340082
rect 259092 338904 259144 338910
rect 259092 338846 259144 338852
rect 259184 335640 259236 335646
rect 259012 335566 259132 335594
rect 259184 335582 259236 335588
rect 259000 335504 259052 335510
rect 259000 335446 259052 335452
rect 258816 328432 258868 328438
rect 258816 328374 258868 328380
rect 258724 326392 258776 326398
rect 258724 326334 258776 326340
rect 258828 322402 258856 328374
rect 258736 322374 258856 322402
rect 258736 317558 258764 322374
rect 258724 317552 258776 317558
rect 258724 317494 258776 317500
rect 258908 317552 258960 317558
rect 258908 317494 258960 317500
rect 258920 315994 258948 317494
rect 258908 315988 258960 315994
rect 258908 315930 258960 315936
rect 258816 298172 258868 298178
rect 258816 298114 258868 298120
rect 258828 298081 258856 298114
rect 258814 298072 258870 298081
rect 258814 298007 258870 298016
rect 258722 297936 258778 297945
rect 258722 297871 258778 297880
rect 258736 293162 258764 297871
rect 258736 293134 258948 293162
rect 258920 287026 258948 293134
rect 258908 287020 258960 287026
rect 258908 286962 258960 286968
rect 258724 277432 258776 277438
rect 258724 277374 258776 277380
rect 258736 258126 258764 277374
rect 258632 258120 258684 258126
rect 258632 258062 258684 258068
rect 258724 258120 258776 258126
rect 258724 258062 258776 258068
rect 258644 249898 258672 258062
rect 258632 249892 258684 249898
rect 258632 249834 258684 249840
rect 258724 249824 258776 249830
rect 258776 249772 258856 249778
rect 258724 249766 258856 249772
rect 258736 249762 258856 249766
rect 258736 249756 258868 249762
rect 258736 249750 258816 249756
rect 258816 249698 258868 249704
rect 258816 240236 258868 240242
rect 258816 240178 258868 240184
rect 258828 240106 258856 240178
rect 258632 240100 258684 240106
rect 258632 240042 258684 240048
rect 258816 240100 258868 240106
rect 258816 240042 258868 240048
rect 258644 230625 258672 240042
rect 258630 230616 258686 230625
rect 258630 230551 258686 230560
rect 258722 230480 258778 230489
rect 258722 230415 258778 230424
rect 258736 202910 258764 230415
rect 258724 202904 258776 202910
rect 258724 202846 258776 202852
rect 258816 202904 258868 202910
rect 258816 202846 258868 202852
rect 258828 191894 258856 202846
rect 258816 191888 258868 191894
rect 258816 191830 258868 191836
rect 258908 191888 258960 191894
rect 258908 191830 258960 191836
rect 258920 186386 258948 191830
rect 258908 186380 258960 186386
rect 258908 186322 258960 186328
rect 258908 186244 258960 186250
rect 258908 186186 258960 186192
rect 258920 172582 258948 186186
rect 258816 172576 258868 172582
rect 258816 172518 258868 172524
rect 258908 172576 258960 172582
rect 258908 172518 258960 172524
rect 258828 164393 258856 172518
rect 258814 164384 258870 164393
rect 258814 164319 258870 164328
rect 258814 164248 258870 164257
rect 258814 164183 258870 164192
rect 258828 157486 258856 164183
rect 258816 157480 258868 157486
rect 258816 157422 258868 157428
rect 258816 157344 258868 157350
rect 258816 157286 258868 157292
rect 258828 143546 258856 157286
rect 258816 143540 258868 143546
rect 258816 143482 258868 143488
rect 258908 138644 258960 138650
rect 258908 138586 258960 138592
rect 258920 125662 258948 138586
rect 258816 125656 258868 125662
rect 258816 125598 258868 125604
rect 258908 125656 258960 125662
rect 258908 125598 258960 125604
rect 258828 120714 258856 125598
rect 258828 120686 258948 120714
rect 258920 115938 258948 120686
rect 258908 115932 258960 115938
rect 258908 115874 258960 115880
rect 258908 106344 258960 106350
rect 258908 106286 258960 106292
rect 258920 103494 258948 106286
rect 258908 103488 258960 103494
rect 258908 103430 258960 103436
rect 258908 93900 258960 93906
rect 258908 93842 258960 93848
rect 258920 93809 258948 93842
rect 258722 93800 258778 93809
rect 258722 93735 258778 93744
rect 258906 93800 258962 93809
rect 258906 93735 258962 93744
rect 258736 84250 258764 93735
rect 258724 84244 258776 84250
rect 258724 84186 258776 84192
rect 258908 84244 258960 84250
rect 258908 84186 258960 84192
rect 258920 76022 258948 84186
rect 258908 76016 258960 76022
rect 258908 75958 258960 75964
rect 258816 75880 258868 75886
rect 258816 75822 258868 75828
rect 258828 64938 258856 75822
rect 258816 64932 258868 64938
rect 258816 64874 258868 64880
rect 258908 64932 258960 64938
rect 258908 64874 258960 64880
rect 258920 60178 258948 64874
rect 258908 60172 258960 60178
rect 258908 60114 258960 60120
rect 258908 60036 258960 60042
rect 258908 59978 258960 59984
rect 258920 37330 258948 59978
rect 258816 37324 258868 37330
rect 258816 37266 258868 37272
rect 258908 37324 258960 37330
rect 258908 37266 258960 37272
rect 258828 6730 258856 37266
rect 258816 6724 258868 6730
rect 258816 6666 258868 6672
rect 258632 5500 258684 5506
rect 258632 5442 258684 5448
rect 257988 5364 258040 5370
rect 257988 5306 258040 5312
rect 257896 5296 257948 5302
rect 257896 5238 257948 5244
rect 258644 480 258672 5442
rect 259012 4418 259040 335446
rect 259104 4554 259132 335566
rect 259092 4548 259144 4554
rect 259092 4490 259144 4496
rect 259000 4412 259052 4418
rect 259000 4354 259052 4360
rect 259196 4350 259224 335582
rect 259288 335442 259316 340054
rect 259460 338700 259512 338706
rect 259460 338642 259512 338648
rect 259276 335436 259328 335442
rect 259276 335378 259328 335384
rect 259368 330744 259420 330750
rect 259368 330686 259420 330692
rect 259276 326392 259328 326398
rect 259276 326334 259328 326340
rect 259288 4962 259316 326334
rect 259276 4956 259328 4962
rect 259276 4898 259328 4904
rect 259184 4344 259236 4350
rect 259184 4286 259236 4292
rect 259380 4214 259408 330686
rect 259472 326466 259500 338642
rect 259644 335640 259696 335646
rect 259644 335582 259696 335588
rect 259460 326460 259512 326466
rect 259460 326402 259512 326408
rect 259656 326210 259684 335582
rect 259748 326398 259776 340054
rect 259840 338706 259868 340068
rect 259932 340054 260130 340082
rect 260208 340054 260314 340082
rect 260392 340054 260590 340082
rect 259828 338700 259880 338706
rect 259828 338642 259880 338648
rect 259736 326392 259788 326398
rect 259932 326380 259960 340054
rect 260208 331294 260236 340054
rect 260392 335646 260420 340054
rect 260380 335640 260432 335646
rect 260380 335582 260432 335588
rect 260196 331288 260248 331294
rect 260196 331230 260248 331236
rect 260012 331220 260064 331226
rect 260012 331162 260064 331168
rect 260024 326618 260052 331162
rect 260024 326590 260696 326618
rect 260564 326460 260616 326466
rect 260564 326402 260616 326408
rect 259932 326352 260512 326380
rect 259736 326334 259788 326340
rect 259656 326182 259776 326210
rect 259748 321570 259776 326182
rect 259736 321564 259788 321570
rect 259736 321506 259788 321512
rect 260380 321564 260432 321570
rect 260380 321506 260432 321512
rect 260392 317422 260420 321506
rect 260380 317416 260432 317422
rect 260380 317358 260432 317364
rect 260380 307828 260432 307834
rect 260380 307770 260432 307776
rect 260392 302138 260420 307770
rect 260300 302110 260420 302138
rect 260300 299470 260328 302110
rect 260288 299464 260340 299470
rect 260288 299406 260340 299412
rect 260380 289876 260432 289882
rect 260380 289818 260432 289824
rect 260392 285002 260420 289818
rect 260300 284974 260420 285002
rect 260300 273290 260328 284974
rect 260288 273284 260340 273290
rect 260288 273226 260340 273232
rect 260380 265328 260432 265334
rect 260380 265270 260432 265276
rect 260392 248441 260420 265270
rect 260194 248432 260250 248441
rect 260194 248367 260250 248376
rect 260378 248432 260434 248441
rect 260378 248367 260434 248376
rect 260208 240310 260236 248367
rect 260196 240304 260248 240310
rect 260196 240246 260248 240252
rect 260288 240168 260340 240174
rect 260288 240110 260340 240116
rect 260300 234682 260328 240110
rect 260208 234654 260328 234682
rect 260208 229226 260236 234654
rect 260196 229220 260248 229226
rect 260196 229162 260248 229168
rect 260380 229220 260432 229226
rect 260380 229162 260432 229168
rect 260392 229090 260420 229162
rect 260380 229084 260432 229090
rect 260380 229026 260432 229032
rect 260380 224256 260432 224262
rect 260380 224198 260432 224204
rect 260392 219434 260420 224198
rect 260380 219428 260432 219434
rect 260380 219370 260432 219376
rect 260380 214532 260432 214538
rect 260380 214474 260432 214480
rect 260392 202910 260420 214474
rect 260288 202904 260340 202910
rect 260288 202846 260340 202852
rect 260380 202904 260432 202910
rect 260380 202846 260432 202852
rect 260300 196738 260328 202846
rect 260208 196710 260328 196738
rect 260208 191826 260236 196710
rect 260196 191820 260248 191826
rect 260196 191762 260248 191768
rect 260288 183524 260340 183530
rect 260288 183466 260340 183472
rect 260300 182170 260328 183466
rect 260288 182164 260340 182170
rect 260288 182106 260340 182112
rect 260288 173868 260340 173874
rect 260288 173810 260340 173816
rect 260300 172530 260328 173810
rect 260300 172502 260420 172530
rect 260392 160070 260420 172502
rect 260380 160064 260432 160070
rect 260380 160006 260432 160012
rect 260288 159996 260340 160002
rect 260288 159938 260340 159944
rect 260300 158710 260328 159938
rect 260288 158704 260340 158710
rect 260288 158646 260340 158652
rect 260288 149116 260340 149122
rect 260288 149058 260340 149064
rect 260300 142186 260328 149058
rect 260288 142180 260340 142186
rect 260288 142122 260340 142128
rect 260288 142044 260340 142050
rect 260288 141986 260340 141992
rect 260300 140842 260328 141986
rect 260208 140814 260328 140842
rect 260208 139398 260236 140814
rect 260196 139392 260248 139398
rect 260196 139334 260248 139340
rect 260288 129804 260340 129810
rect 260288 129746 260340 129752
rect 260300 120714 260328 129746
rect 260300 120686 260420 120714
rect 260392 115938 260420 120686
rect 260380 115932 260432 115938
rect 260380 115874 260432 115880
rect 260380 106344 260432 106350
rect 260380 106286 260432 106292
rect 260392 100042 260420 106286
rect 260300 100014 260420 100042
rect 259458 87000 259514 87009
rect 259458 86935 259514 86944
rect 259472 86873 259500 86935
rect 259458 86864 259514 86873
rect 259458 86799 259514 86808
rect 260300 85610 260328 100014
rect 260288 85604 260340 85610
rect 260288 85546 260340 85552
rect 260380 85604 260432 85610
rect 260380 85546 260432 85552
rect 260392 76022 260420 85546
rect 260380 76016 260432 76022
rect 260380 75958 260432 75964
rect 260288 75880 260340 75886
rect 260288 75822 260340 75828
rect 260300 66366 260328 75822
rect 260288 66360 260340 66366
rect 260288 66302 260340 66308
rect 260196 66292 260248 66298
rect 260196 66234 260248 66240
rect 260208 64870 260236 66234
rect 260196 64864 260248 64870
rect 260196 64806 260248 64812
rect 260380 64864 260432 64870
rect 260380 64806 260432 64812
rect 259458 40216 259514 40225
rect 259458 40151 259514 40160
rect 259472 40089 259500 40151
rect 259458 40080 259514 40089
rect 259458 40015 259514 40024
rect 259458 17096 259514 17105
rect 259458 17031 259514 17040
rect 259472 16697 259500 17031
rect 259458 16688 259514 16697
rect 259458 16623 259514 16632
rect 260392 6526 260420 64806
rect 260484 6662 260512 326352
rect 260576 6798 260604 326402
rect 260564 6792 260616 6798
rect 260564 6734 260616 6740
rect 260472 6656 260524 6662
rect 260472 6598 260524 6604
rect 260380 6520 260432 6526
rect 260380 6462 260432 6468
rect 259828 5432 259880 5438
rect 259828 5374 259880 5380
rect 259368 4208 259420 4214
rect 259368 4150 259420 4156
rect 259840 480 259868 5374
rect 260668 4758 260696 326590
rect 260852 326466 260880 340068
rect 260944 340054 261050 340082
rect 260840 326460 260892 326466
rect 260840 326402 260892 326408
rect 260748 326392 260800 326398
rect 260748 326334 260800 326340
rect 260760 5030 260788 326334
rect 260944 326330 260972 340054
rect 261312 335850 261340 340068
rect 261404 340054 261602 340082
rect 261680 340054 261786 340082
rect 261864 340054 262062 340082
rect 262338 340054 262444 340082
rect 261300 335844 261352 335850
rect 261300 335786 261352 335792
rect 261300 335708 261352 335714
rect 261300 335650 261352 335656
rect 261208 335640 261260 335646
rect 261208 335582 261260 335588
rect 261116 333328 261168 333334
rect 261116 333270 261168 333276
rect 260932 326324 260984 326330
rect 260932 326266 260984 326272
rect 261128 324494 261156 333270
rect 261220 326398 261248 335582
rect 261208 326392 261260 326398
rect 261312 326380 261340 335650
rect 261404 333334 261432 340054
rect 261680 335646 261708 340054
rect 261668 335640 261720 335646
rect 261668 335582 261720 335588
rect 261392 333328 261444 333334
rect 261392 333270 261444 333276
rect 261864 333198 261892 340054
rect 262220 335708 262272 335714
rect 262220 335650 262272 335656
rect 261392 333192 261444 333198
rect 261392 333134 261444 333140
rect 261852 333192 261904 333198
rect 261852 333134 261904 333140
rect 261404 326618 261432 333134
rect 261404 326590 261984 326618
rect 261852 326460 261904 326466
rect 261852 326402 261904 326408
rect 261312 326352 261800 326380
rect 261208 326334 261260 326340
rect 261116 324488 261168 324494
rect 261116 324430 261168 324436
rect 261576 324488 261628 324494
rect 261576 324430 261628 324436
rect 261588 318866 261616 324430
rect 261588 318838 261708 318866
rect 261680 317422 261708 318838
rect 261668 317416 261720 317422
rect 261668 317358 261720 317364
rect 261576 299532 261628 299538
rect 261576 299474 261628 299480
rect 261588 294794 261616 299474
rect 261496 294766 261616 294794
rect 261496 289814 261524 294766
rect 261484 289808 261536 289814
rect 261484 289750 261536 289756
rect 261576 289808 261628 289814
rect 261576 289750 261628 289756
rect 261588 278769 261616 289750
rect 261390 278760 261446 278769
rect 261390 278695 261446 278704
rect 261574 278760 261630 278769
rect 261574 278695 261630 278704
rect 261404 269142 261432 278695
rect 261392 269136 261444 269142
rect 261392 269078 261444 269084
rect 261668 269136 261720 269142
rect 261668 269078 261720 269084
rect 261680 265554 261708 269078
rect 261588 265526 261708 265554
rect 261588 254810 261616 265526
rect 261496 254782 261616 254810
rect 261496 240174 261524 254782
rect 261484 240168 261536 240174
rect 261484 240110 261536 240116
rect 261576 240168 261628 240174
rect 261576 240110 261628 240116
rect 261588 238746 261616 240110
rect 261576 238740 261628 238746
rect 261576 238682 261628 238688
rect 261576 234592 261628 234598
rect 261576 234534 261628 234540
rect 261588 229106 261616 234534
rect 261588 229078 261708 229106
rect 261680 227066 261708 229078
rect 261588 227038 261708 227066
rect 261588 219434 261616 227038
rect 261576 219428 261628 219434
rect 261576 219370 261628 219376
rect 261576 215280 261628 215286
rect 261576 215222 261628 215228
rect 261588 209794 261616 215222
rect 261588 209766 261708 209794
rect 261680 203658 261708 209766
rect 261576 203652 261628 203658
rect 261576 203594 261628 203600
rect 261668 203652 261720 203658
rect 261668 203594 261720 203600
rect 261588 196738 261616 203594
rect 261496 196710 261616 196738
rect 261496 190466 261524 196710
rect 261484 190460 261536 190466
rect 261484 190402 261536 190408
rect 261484 182164 261536 182170
rect 261484 182106 261536 182112
rect 261496 180826 261524 182106
rect 261496 180798 261616 180826
rect 261588 175930 261616 180798
rect 261588 175902 261708 175930
rect 261680 164354 261708 175902
rect 261668 164348 261720 164354
rect 261668 164290 261720 164296
rect 261576 164280 261628 164286
rect 261576 164222 261628 164228
rect 261588 162858 261616 164222
rect 261576 162852 261628 162858
rect 261576 162794 261628 162800
rect 261668 162852 261720 162858
rect 261668 162794 261720 162800
rect 261680 142202 261708 162794
rect 261588 142174 261708 142202
rect 261588 131238 261616 142174
rect 261484 131232 261536 131238
rect 261484 131174 261536 131180
rect 261576 131232 261628 131238
rect 261576 131174 261628 131180
rect 261496 131102 261524 131174
rect 261484 131096 261536 131102
rect 261484 131038 261536 131044
rect 261484 122732 261536 122738
rect 261484 122674 261536 122680
rect 261496 121446 261524 122674
rect 261484 121440 261536 121446
rect 261484 121382 261536 121388
rect 261484 111852 261536 111858
rect 261484 111794 261536 111800
rect 261496 103630 261524 111794
rect 261484 103624 261536 103630
rect 261484 103566 261536 103572
rect 261392 103556 261444 103562
rect 261392 103498 261444 103504
rect 261404 99822 261432 103498
rect 261392 99816 261444 99822
rect 261392 99758 261444 99764
rect 261668 85536 261720 85542
rect 261668 85478 261720 85484
rect 261680 84182 261708 85478
rect 261668 84176 261720 84182
rect 261668 84118 261720 84124
rect 261668 74656 261720 74662
rect 261668 74598 261720 74604
rect 261680 56030 261708 74598
rect 261668 56024 261720 56030
rect 261668 55966 261720 55972
rect 261576 46980 261628 46986
rect 261576 46922 261628 46928
rect 261588 42158 261616 46922
rect 261576 42152 261628 42158
rect 261576 42094 261628 42100
rect 261668 35964 261720 35970
rect 261668 35906 261720 35912
rect 261680 6390 261708 35906
rect 261772 6458 261800 326352
rect 261864 6594 261892 326402
rect 261852 6588 261904 6594
rect 261852 6530 261904 6536
rect 261760 6452 261812 6458
rect 261760 6394 261812 6400
rect 261668 6384 261720 6390
rect 261668 6326 261720 6332
rect 261956 6322 261984 326590
rect 262036 326392 262088 326398
rect 262036 326334 262088 326340
rect 261944 6316 261996 6322
rect 261944 6258 261996 6264
rect 261024 5364 261076 5370
rect 261024 5306 261076 5312
rect 260748 5024 260800 5030
rect 260748 4966 260800 4972
rect 260656 4752 260708 4758
rect 260656 4694 260708 4700
rect 261036 480 261064 5306
rect 262048 4826 262076 326334
rect 262232 326330 262260 335650
rect 262416 335646 262444 340054
rect 262404 335640 262456 335646
rect 262404 335582 262456 335588
rect 262404 335504 262456 335510
rect 262404 335446 262456 335452
rect 262416 326534 262444 335446
rect 262404 326528 262456 326534
rect 262404 326470 262456 326476
rect 262128 326324 262180 326330
rect 262128 326266 262180 326272
rect 262220 326324 262272 326330
rect 262220 326266 262272 326272
rect 262140 4894 262168 326266
rect 262508 326262 262536 340068
rect 262588 339108 262640 339114
rect 262588 339050 262640 339056
rect 262600 326466 262628 339050
rect 262968 336977 262996 340190
rect 279528 340190 279726 340218
rect 282472 340202 282670 340218
rect 300596 340202 300794 340218
rect 281724 340196 281776 340202
rect 263060 339114 263088 340068
rect 263152 340054 263258 340082
rect 263336 340054 263534 340082
rect 263612 340054 263810 340082
rect 263048 339108 263100 339114
rect 263048 339050 263100 339056
rect 262954 336968 263010 336977
rect 262954 336903 263010 336912
rect 262770 336832 262826 336841
rect 262770 336767 262826 336776
rect 262680 335640 262732 335646
rect 262680 335582 262732 335588
rect 262588 326460 262640 326466
rect 262588 326402 262640 326408
rect 262692 326398 262720 335582
rect 262784 333742 262812 336767
rect 263152 335510 263180 340054
rect 263336 335714 263364 340054
rect 263324 335708 263376 335714
rect 263324 335650 263376 335656
rect 263140 335504 263192 335510
rect 263140 335446 263192 335452
rect 262772 333736 262824 333742
rect 262772 333678 262824 333684
rect 263324 326528 263376 326534
rect 263324 326470 263376 326476
rect 262680 326392 262732 326398
rect 262680 326334 262732 326340
rect 263232 326392 263284 326398
rect 263232 326334 263284 326340
rect 263140 326324 263192 326330
rect 263140 326266 263192 326272
rect 262496 326256 262548 326262
rect 262496 326198 262548 326204
rect 262864 325712 262916 325718
rect 262864 325654 262916 325660
rect 262876 322250 262904 325654
rect 262864 322244 262916 322250
rect 262864 322186 262916 322192
rect 263048 322244 263100 322250
rect 263048 322186 263100 322192
rect 263060 263650 263088 322186
rect 262968 263622 263088 263650
rect 262968 263514 262996 263622
rect 262968 263486 263088 263514
rect 263060 244338 263088 263486
rect 262968 244310 263088 244338
rect 262968 244202 262996 244310
rect 262968 244174 263088 244202
rect 263060 225026 263088 244174
rect 262968 224998 263088 225026
rect 262968 224890 262996 224998
rect 262968 224862 263088 224890
rect 263060 205630 263088 224862
rect 262864 205624 262916 205630
rect 262864 205566 262916 205572
rect 263048 205624 263100 205630
rect 263048 205566 263100 205572
rect 262876 200161 262904 205566
rect 262862 200152 262918 200161
rect 262862 200087 262918 200096
rect 263046 200152 263102 200161
rect 263046 200087 263102 200096
rect 263060 190466 263088 200087
rect 263048 190460 263100 190466
rect 263048 190402 263100 190408
rect 263048 180872 263100 180878
rect 263048 180814 263100 180820
rect 263060 118046 263088 180814
rect 263048 118040 263100 118046
rect 263048 117982 263100 117988
rect 263048 104916 263100 104922
rect 263048 104858 263100 104864
rect 263060 103494 263088 104858
rect 263048 103488 263100 103494
rect 263048 103430 263100 103436
rect 263048 93900 263100 93906
rect 263048 93842 263100 93848
rect 263060 89826 263088 93842
rect 263048 89820 263100 89826
rect 263048 89762 263100 89768
rect 263048 89684 263100 89690
rect 263048 89626 263100 89632
rect 263060 83026 263088 89626
rect 263048 83020 263100 83026
rect 263048 82962 263100 82968
rect 263048 67652 263100 67658
rect 263048 67594 263100 67600
rect 263060 41426 263088 67594
rect 262968 41398 263088 41426
rect 262968 31822 262996 41398
rect 262956 31816 263008 31822
rect 262956 31758 263008 31764
rect 263048 31680 263100 31686
rect 263048 31622 263100 31628
rect 263060 24154 263088 31622
rect 262968 24126 263088 24154
rect 262968 6254 262996 24126
rect 262956 6248 263008 6254
rect 262956 6190 263008 6196
rect 263152 6186 263180 326266
rect 263140 6180 263192 6186
rect 263140 6122 263192 6128
rect 262220 5296 262272 5302
rect 262220 5238 262272 5244
rect 262128 4888 262180 4894
rect 262128 4830 262180 4836
rect 262036 4820 262088 4826
rect 262036 4762 262088 4768
rect 262232 480 262260 5238
rect 263244 4486 263272 326334
rect 263336 4622 263364 326470
rect 263416 326460 263468 326466
rect 263416 326402 263468 326408
rect 263428 4690 263456 326402
rect 263612 326398 263640 340054
rect 263980 335646 264008 340068
rect 264072 340054 264270 340082
rect 264546 340054 264652 340082
rect 263968 335640 264020 335646
rect 263968 335582 264020 335588
rect 264072 333282 264100 340054
rect 263704 333254 264100 333282
rect 263704 328438 263732 333254
rect 263876 332376 263928 332382
rect 263876 332318 263928 332324
rect 263692 328432 263744 328438
rect 263692 328374 263744 328380
rect 263784 328364 263836 328370
rect 263784 328306 263836 328312
rect 263600 326392 263652 326398
rect 263600 326334 263652 326340
rect 263508 326256 263560 326262
rect 263508 326198 263560 326204
rect 263416 4684 263468 4690
rect 263416 4626 263468 4632
rect 263324 4616 263376 4622
rect 263324 4558 263376 4564
rect 263520 4554 263548 326198
rect 263796 313546 263824 328306
rect 263888 326346 263916 332318
rect 264624 332194 264652 340054
rect 264716 332382 264744 340068
rect 264888 335640 264940 335646
rect 264888 335582 264940 335588
rect 264704 332376 264756 332382
rect 264704 332318 264756 332324
rect 264624 332166 264744 332194
rect 263888 326318 264560 326346
rect 264532 316690 264560 326318
rect 264532 316662 264652 316690
rect 263784 313540 263836 313546
rect 263784 313482 263836 313488
rect 264520 313540 264572 313546
rect 264520 313482 264572 313488
rect 264532 307766 264560 313482
rect 264520 307760 264572 307766
rect 264520 307702 264572 307708
rect 264520 298172 264572 298178
rect 264520 298114 264572 298120
rect 264532 278730 264560 298114
rect 264520 278724 264572 278730
rect 264520 278666 264572 278672
rect 264520 269136 264572 269142
rect 264334 269104 264390 269113
rect 264334 269039 264390 269048
rect 264518 269104 264520 269113
rect 264572 269104 264574 269113
rect 264518 269039 264574 269048
rect 264348 259486 264376 269039
rect 264336 259480 264388 259486
rect 264336 259422 264388 259428
rect 264520 259480 264572 259486
rect 264520 259422 264572 259428
rect 264532 249801 264560 259422
rect 264334 249792 264390 249801
rect 264334 249727 264390 249736
rect 264518 249792 264574 249801
rect 264518 249727 264574 249736
rect 264348 240174 264376 249727
rect 264336 240168 264388 240174
rect 264336 240110 264388 240116
rect 264520 240168 264572 240174
rect 264520 240110 264572 240116
rect 264532 211138 264560 240110
rect 264336 211132 264388 211138
rect 264336 211074 264388 211080
rect 264520 211132 264572 211138
rect 264520 211074 264572 211080
rect 264348 201521 264376 211074
rect 264334 201512 264390 201521
rect 264334 201447 264336 201456
rect 264388 201447 264390 201456
rect 264518 201512 264574 201521
rect 264518 201447 264520 201456
rect 264336 201418 264388 201424
rect 264572 201447 264574 201456
rect 264520 201418 264572 201424
rect 264348 191865 264376 201418
rect 264334 191856 264390 191865
rect 264334 191791 264336 191800
rect 264388 191791 264390 191800
rect 264518 191856 264574 191865
rect 264518 191791 264520 191800
rect 264336 191762 264388 191768
rect 264572 191791 264574 191800
rect 264520 191762 264572 191768
rect 264348 182209 264376 191762
rect 264334 182200 264390 182209
rect 264334 182135 264390 182144
rect 264518 182200 264574 182209
rect 264518 182135 264574 182144
rect 264532 180810 264560 182135
rect 264520 180804 264572 180810
rect 264520 180746 264572 180752
rect 264520 171148 264572 171154
rect 264520 171090 264572 171096
rect 264532 151774 264560 171090
rect 264520 151768 264572 151774
rect 264520 151710 264572 151716
rect 264520 142180 264572 142186
rect 264520 142122 264572 142128
rect 264532 122806 264560 142122
rect 264520 122800 264572 122806
rect 264520 122742 264572 122748
rect 264520 113212 264572 113218
rect 264520 113154 264572 113160
rect 264532 103494 264560 113154
rect 264520 103488 264572 103494
rect 264520 103430 264572 103436
rect 264428 93900 264480 93906
rect 264428 93842 264480 93848
rect 264440 85610 264468 93842
rect 264428 85604 264480 85610
rect 264428 85546 264480 85552
rect 264520 85604 264572 85610
rect 264520 85546 264572 85552
rect 264532 84182 264560 85546
rect 264520 84176 264572 84182
rect 264520 84118 264572 84124
rect 264520 74588 264572 74594
rect 264520 74530 264572 74536
rect 264532 64870 264560 74530
rect 264520 64864 264572 64870
rect 264520 64806 264572 64812
rect 264520 46980 264572 46986
rect 264520 46922 264572 46928
rect 264532 45558 264560 46922
rect 264520 45552 264572 45558
rect 264520 45494 264572 45500
rect 264428 35964 264480 35970
rect 264428 35906 264480 35912
rect 264440 29034 264468 35906
rect 264428 29028 264480 29034
rect 264428 28970 264480 28976
rect 264520 29028 264572 29034
rect 264520 28970 264572 28976
rect 264242 16280 264298 16289
rect 264242 16215 264298 16224
rect 264256 15609 264284 16215
rect 264242 15600 264298 15609
rect 264242 15535 264298 15544
rect 264532 7954 264560 28970
rect 264520 7948 264572 7954
rect 264520 7890 264572 7896
rect 264624 5370 264652 316662
rect 264716 5438 264744 332166
rect 264796 326392 264848 326398
rect 264796 326334 264848 326340
rect 264704 5432 264756 5438
rect 264704 5374 264756 5380
rect 264612 5364 264664 5370
rect 264612 5306 264664 5312
rect 263508 4548 263560 4554
rect 263508 4490 263560 4496
rect 263232 4480 263284 4486
rect 263232 4422 263284 4428
rect 263324 4412 263376 4418
rect 263324 4354 263376 4360
rect 263336 3074 263364 4354
rect 264808 4214 264836 326334
rect 264900 5506 264928 335582
rect 264992 326466 265020 340068
rect 265164 335640 265216 335646
rect 265164 335582 265216 335588
rect 265072 335028 265124 335034
rect 265072 334970 265124 334976
rect 264980 326460 265032 326466
rect 264980 326402 265032 326408
rect 265084 326398 265112 334970
rect 265072 326392 265124 326398
rect 265072 326334 265124 326340
rect 265176 326330 265204 335582
rect 265268 328234 265296 340068
rect 265360 340054 265466 340082
rect 265544 340054 265742 340082
rect 266018 340054 266124 340082
rect 265360 335646 265388 340054
rect 265348 335640 265400 335646
rect 265348 335582 265400 335588
rect 265544 328506 265572 340054
rect 266096 333418 266124 340054
rect 266188 335034 266216 340068
rect 266372 340054 266478 340082
rect 266556 340054 266754 340082
rect 266832 340054 266938 340082
rect 267214 340054 267320 340082
rect 266372 338201 266400 340054
rect 266358 338192 266414 338201
rect 266358 338127 266414 338136
rect 266360 335640 266412 335646
rect 266360 335582 266412 335588
rect 266176 335028 266228 335034
rect 266176 334970 266228 334976
rect 266096 333390 266308 333418
rect 265440 328500 265492 328506
rect 265440 328442 265492 328448
rect 265532 328500 265584 328506
rect 265532 328442 265584 328448
rect 265452 328386 265480 328442
rect 265452 328358 265664 328386
rect 265256 328228 265308 328234
rect 265256 328170 265308 328176
rect 265164 326324 265216 326330
rect 265164 326266 265216 326272
rect 265636 318850 265664 328358
rect 266084 328228 266136 328234
rect 266084 328170 266136 328176
rect 265900 326460 265952 326466
rect 265900 326402 265952 326408
rect 265624 318844 265676 318850
rect 265624 318786 265676 318792
rect 265808 318708 265860 318714
rect 265808 318650 265860 318656
rect 265820 317422 265848 318650
rect 265808 317416 265860 317422
rect 265808 317358 265860 317364
rect 265808 307896 265860 307902
rect 265808 307838 265860 307844
rect 265820 307766 265848 307838
rect 265808 307760 265860 307766
rect 265808 307702 265860 307708
rect 265808 298172 265860 298178
rect 265808 298114 265860 298120
rect 265820 288386 265848 298114
rect 265808 288380 265860 288386
rect 265808 288322 265860 288328
rect 265808 278860 265860 278866
rect 265808 278802 265860 278808
rect 265820 278730 265848 278802
rect 265808 278724 265860 278730
rect 265808 278666 265860 278672
rect 265808 269136 265860 269142
rect 265622 269104 265678 269113
rect 265622 269039 265678 269048
rect 265806 269104 265808 269113
rect 265860 269104 265862 269113
rect 265806 269039 265862 269048
rect 265636 259486 265664 269039
rect 265624 259480 265676 259486
rect 265624 259422 265676 259428
rect 265808 259480 265860 259486
rect 265808 259422 265860 259428
rect 265820 253230 265848 259422
rect 265624 253224 265676 253230
rect 265624 253166 265676 253172
rect 265808 253224 265860 253230
rect 265808 253166 265860 253172
rect 265636 248441 265664 253166
rect 265622 248432 265678 248441
rect 265622 248367 265678 248376
rect 265806 248432 265862 248441
rect 265806 248367 265862 248376
rect 265820 238746 265848 248367
rect 265624 238740 265676 238746
rect 265624 238682 265676 238688
rect 265808 238740 265860 238746
rect 265808 238682 265860 238688
rect 265636 229129 265664 238682
rect 265622 229120 265678 229129
rect 265622 229055 265678 229064
rect 265806 229120 265862 229129
rect 265806 229055 265862 229064
rect 265820 219434 265848 229055
rect 265624 219428 265676 219434
rect 265624 219370 265676 219376
rect 265808 219428 265860 219434
rect 265808 219370 265860 219376
rect 265636 209817 265664 219370
rect 265622 209808 265678 209817
rect 265622 209743 265678 209752
rect 265806 209808 265862 209817
rect 265806 209743 265862 209752
rect 265820 191826 265848 209743
rect 265624 191820 265676 191826
rect 265624 191762 265676 191768
rect 265808 191820 265860 191826
rect 265808 191762 265860 191768
rect 265636 182209 265664 191762
rect 265622 182200 265678 182209
rect 265622 182135 265678 182144
rect 265806 182200 265862 182209
rect 265806 182135 265862 182144
rect 265820 180810 265848 182135
rect 265808 180804 265860 180810
rect 265808 180746 265860 180752
rect 265808 171148 265860 171154
rect 265808 171090 265860 171096
rect 265820 122806 265848 171090
rect 265808 122800 265860 122806
rect 265808 122742 265860 122748
rect 265808 113212 265860 113218
rect 265808 113154 265860 113160
rect 265820 103494 265848 113154
rect 265808 103488 265860 103494
rect 265808 103430 265860 103436
rect 265716 95192 265768 95198
rect 265716 95134 265768 95140
rect 265728 85610 265756 95134
rect 265716 85604 265768 85610
rect 265716 85546 265768 85552
rect 265808 85604 265860 85610
rect 265808 85546 265860 85552
rect 265820 84182 265848 85546
rect 265808 84176 265860 84182
rect 265808 84118 265860 84124
rect 265806 74624 265862 74633
rect 265806 74559 265862 74568
rect 265820 74526 265848 74559
rect 265624 74520 265676 74526
rect 265624 74462 265676 74468
rect 265808 74520 265860 74526
rect 265808 74462 265860 74468
rect 265636 64977 265664 74462
rect 265622 64968 265678 64977
rect 265622 64903 265678 64912
rect 265806 64968 265862 64977
rect 265806 64903 265862 64912
rect 265820 64870 265848 64903
rect 265808 64864 265860 64870
rect 265808 64806 265860 64812
rect 265808 55344 265860 55350
rect 265808 55286 265860 55292
rect 265820 55214 265848 55286
rect 265808 55208 265860 55214
rect 265808 55150 265860 55156
rect 265808 45620 265860 45626
rect 265808 45562 265860 45568
rect 265820 37398 265848 45562
rect 265808 37392 265860 37398
rect 265808 37334 265860 37340
rect 265716 35964 265768 35970
rect 265716 35906 265768 35912
rect 265728 29034 265756 35906
rect 265716 29028 265768 29034
rect 265716 28970 265768 28976
rect 265808 29028 265860 29034
rect 265808 28970 265860 28976
rect 265820 7818 265848 28970
rect 265912 7886 265940 326402
rect 265992 326392 266044 326398
rect 265992 326334 266044 326340
rect 265900 7880 265952 7886
rect 265900 7822 265952 7828
rect 265808 7812 265860 7818
rect 265808 7754 265860 7760
rect 264888 5500 264940 5506
rect 264888 5442 264940 5448
rect 266004 4826 266032 326334
rect 266096 5302 266124 328170
rect 266176 326324 266228 326330
rect 266176 326266 266228 326272
rect 266084 5296 266136 5302
rect 266084 5238 266136 5244
rect 266188 5234 266216 326266
rect 266176 5228 266228 5234
rect 266176 5170 266228 5176
rect 266280 5166 266308 333390
rect 266372 326466 266400 335582
rect 266360 326460 266412 326466
rect 266360 326402 266412 326408
rect 266556 326330 266584 340054
rect 266636 335708 266688 335714
rect 266636 335650 266688 335656
rect 266648 326398 266676 335650
rect 266832 335646 266860 340054
rect 266820 335640 266872 335646
rect 266820 335582 266872 335588
rect 266820 335504 266872 335510
rect 266820 335446 266872 335452
rect 266832 327146 266860 335446
rect 266910 328400 266966 328409
rect 266910 328335 266966 328344
rect 266820 327140 266872 327146
rect 266820 327082 266872 327088
rect 266636 326392 266688 326398
rect 266636 326334 266688 326340
rect 266544 326324 266596 326330
rect 266544 326266 266596 326272
rect 266924 321502 266952 328335
rect 266912 321496 266964 321502
rect 266912 321438 266964 321444
rect 267188 321496 267240 321502
rect 267188 321438 267240 321444
rect 267200 304366 267228 321438
rect 267188 304360 267240 304366
rect 267188 304302 267240 304308
rect 267188 304224 267240 304230
rect 267188 304166 267240 304172
rect 267200 227118 267228 304166
rect 267188 227112 267240 227118
rect 267188 227054 267240 227060
rect 267188 226976 267240 226982
rect 267188 226918 267240 226924
rect 267200 207806 267228 226918
rect 267188 207800 267240 207806
rect 267188 207742 267240 207748
rect 267188 207664 267240 207670
rect 267188 207606 267240 207612
rect 266360 84176 266412 84182
rect 266360 84118 266412 84124
rect 266372 74633 266400 84118
rect 266358 74624 266414 74633
rect 266358 74559 266414 74568
rect 267200 38604 267228 207606
rect 267108 38576 267228 38604
rect 267108 29034 267136 38576
rect 267096 29028 267148 29034
rect 267096 28970 267148 28976
rect 267188 29028 267240 29034
rect 267188 28970 267240 28976
rect 267200 19258 267228 28970
rect 267108 19230 267228 19258
rect 267108 9722 267136 19230
rect 267096 9716 267148 9722
rect 267096 9658 267148 9664
rect 267188 9716 267240 9722
rect 267188 9658 267240 9664
rect 267200 7750 267228 9658
rect 267188 7744 267240 7750
rect 267188 7686 267240 7692
rect 267292 7682 267320 340054
rect 267384 340054 267490 340082
rect 267568 340054 267674 340082
rect 267950 340054 268056 340082
rect 267384 335510 267412 340054
rect 267568 335714 267596 340054
rect 267740 338972 267792 338978
rect 267740 338914 267792 338920
rect 267556 335708 267608 335714
rect 267556 335650 267608 335656
rect 267372 335504 267424 335510
rect 267372 335446 267424 335452
rect 267464 327140 267516 327146
rect 267464 327082 267516 327088
rect 267372 326460 267424 326466
rect 267372 326402 267424 326408
rect 267280 7676 267332 7682
rect 267280 7618 267332 7624
rect 267384 5370 267412 326402
rect 267372 5364 267424 5370
rect 267372 5306 267424 5312
rect 266268 5160 266320 5166
rect 266268 5102 266320 5108
rect 267476 4894 267504 327082
rect 267752 326466 267780 338914
rect 267832 335708 267884 335714
rect 267832 335650 267884 335656
rect 267844 327350 267872 335650
rect 267832 327344 267884 327350
rect 267832 327286 267884 327292
rect 267740 326460 267792 326466
rect 267740 326402 267792 326408
rect 268028 326398 268056 340054
rect 268212 338978 268240 340068
rect 268200 338972 268252 338978
rect 268200 338914 268252 338920
rect 268396 335646 268424 340068
rect 268488 340054 268686 340082
rect 268764 340054 268962 340082
rect 269146 340054 269344 340082
rect 268384 335640 268436 335646
rect 268384 335582 268436 335588
rect 268488 333282 268516 340054
rect 268764 335714 268792 340054
rect 269212 335844 269264 335850
rect 269212 335786 269264 335792
rect 268752 335708 268804 335714
rect 268752 335650 268804 335656
rect 269028 335640 269080 335646
rect 269028 335582 269080 335588
rect 268120 333254 268516 333282
rect 267556 326392 267608 326398
rect 267556 326334 267608 326340
rect 268016 326392 268068 326398
rect 268016 326334 268068 326340
rect 267568 5545 267596 326334
rect 267648 326324 267700 326330
rect 267648 326266 267700 326272
rect 267554 5536 267610 5545
rect 267554 5471 267610 5480
rect 267660 5098 267688 326266
rect 268120 324766 268148 333254
rect 268844 327344 268896 327350
rect 268844 327286 268896 327292
rect 268752 326392 268804 326398
rect 268752 326334 268804 326340
rect 268108 324760 268160 324766
rect 268108 324702 268160 324708
rect 268660 324760 268712 324766
rect 268660 324702 268712 324708
rect 268672 304366 268700 324702
rect 268660 304360 268712 304366
rect 268660 304302 268712 304308
rect 268660 304224 268712 304230
rect 268660 304166 268712 304172
rect 268672 227118 268700 304166
rect 268660 227112 268712 227118
rect 268660 227054 268712 227060
rect 268660 226976 268712 226982
rect 268660 226918 268712 226924
rect 268672 207806 268700 226918
rect 268660 207800 268712 207806
rect 268660 207742 268712 207748
rect 268660 207664 268712 207670
rect 268660 207606 268712 207612
rect 267738 63608 267794 63617
rect 267738 63543 267794 63552
rect 267752 63209 267780 63543
rect 267738 63200 267794 63209
rect 267738 63135 267794 63144
rect 267738 40488 267794 40497
rect 267738 40423 267794 40432
rect 267752 40089 267780 40423
rect 267738 40080 267794 40089
rect 267738 40015 267794 40024
rect 268672 38604 268700 207606
rect 268580 38576 268700 38604
rect 268580 29034 268608 38576
rect 268568 29028 268620 29034
rect 268568 28970 268620 28976
rect 268660 29028 268712 29034
rect 268660 28970 268712 28976
rect 268672 19258 268700 28970
rect 268580 19230 268700 19258
rect 268580 9722 268608 19230
rect 268764 16726 268792 326334
rect 268752 16720 268804 16726
rect 268752 16662 268804 16668
rect 268856 16658 268884 327286
rect 268936 326460 268988 326466
rect 268936 326402 268988 326408
rect 268948 16726 268976 326402
rect 268936 16720 268988 16726
rect 268936 16662 268988 16668
rect 269040 16658 269068 335582
rect 269224 326466 269252 335786
rect 269316 335714 269344 340054
rect 269304 335708 269356 335714
rect 269304 335650 269356 335656
rect 269408 335628 269436 340068
rect 269684 335646 269712 340068
rect 269776 340054 269882 340082
rect 269960 340054 270158 340082
rect 270236 340054 270434 340082
rect 269672 335640 269724 335646
rect 269408 335600 269620 335628
rect 269592 327962 269620 335600
rect 269672 335582 269724 335588
rect 269776 335238 269804 340054
rect 269764 335232 269816 335238
rect 269764 335174 269816 335180
rect 269580 327956 269632 327962
rect 269580 327898 269632 327904
rect 269212 326460 269264 326466
rect 269212 326402 269264 326408
rect 268844 16652 268896 16658
rect 268844 16594 268896 16600
rect 269028 16652 269080 16658
rect 269028 16594 269080 16600
rect 268658 16416 268714 16425
rect 269026 16416 269082 16425
rect 268714 16374 269026 16402
rect 268658 16351 268714 16360
rect 269026 16351 269082 16360
rect 268936 13184 268988 13190
rect 268936 13126 268988 13132
rect 268752 13116 268804 13122
rect 268752 13058 268804 13064
rect 268568 9716 268620 9722
rect 268568 9658 268620 9664
rect 268660 9716 268712 9722
rect 268660 9658 268712 9664
rect 268672 9178 268700 9658
rect 268660 9172 268712 9178
rect 268660 9114 268712 9120
rect 268764 7614 268792 13058
rect 268844 12572 268896 12578
rect 268844 12514 268896 12520
rect 268752 7608 268804 7614
rect 268752 7550 268804 7556
rect 268856 5137 268884 12514
rect 268842 5128 268898 5137
rect 267648 5092 267700 5098
rect 268842 5063 268898 5072
rect 267648 5034 267700 5040
rect 268108 4956 268160 4962
rect 268108 4898 268160 4904
rect 267464 4888 267516 4894
rect 267464 4830 267516 4836
rect 265992 4820 266044 4826
rect 265992 4762 266044 4768
rect 265808 4344 265860 4350
rect 265808 4286 265860 4292
rect 264612 4208 264664 4214
rect 264612 4150 264664 4156
rect 264796 4208 264848 4214
rect 264796 4150 264848 4156
rect 263692 3868 263744 3874
rect 263692 3810 263744 3816
rect 263416 3664 263468 3670
rect 263416 3606 263468 3612
rect 263428 3233 263456 3606
rect 263704 3233 263732 3810
rect 263414 3224 263470 3233
rect 263414 3159 263470 3168
rect 263690 3224 263746 3233
rect 263690 3159 263746 3168
rect 263336 3046 263456 3074
rect 263428 480 263456 3046
rect 264624 480 264652 4150
rect 265820 480 265848 4286
rect 267004 4276 267056 4282
rect 267004 4218 267056 4224
rect 267016 480 267044 4218
rect 268120 480 268148 4898
rect 268948 4826 268976 13126
rect 269028 13116 269080 13122
rect 269028 13058 269080 13064
rect 269040 5409 269068 13058
rect 269960 8974 269988 340054
rect 270236 335850 270264 340054
rect 270224 335844 270276 335850
rect 270224 335786 270276 335792
rect 270224 335708 270276 335714
rect 270224 335650 270276 335656
rect 270132 335232 270184 335238
rect 270132 335174 270184 335180
rect 270040 327956 270092 327962
rect 270040 327898 270092 327904
rect 270052 9110 270080 327898
rect 270040 9104 270092 9110
rect 270040 9046 270092 9052
rect 269948 8968 270000 8974
rect 269948 8910 270000 8916
rect 270144 7002 270172 335174
rect 270132 6996 270184 7002
rect 270132 6938 270184 6944
rect 269304 6724 269356 6730
rect 269304 6666 269356 6672
rect 269026 5400 269082 5409
rect 269026 5335 269082 5344
rect 268936 4820 268988 4826
rect 268936 4762 268988 4768
rect 269316 480 269344 6666
rect 270236 5273 270264 335650
rect 270408 335640 270460 335646
rect 270408 335582 270460 335588
rect 270500 335640 270552 335646
rect 270500 335582 270552 335588
rect 270316 326460 270368 326466
rect 270316 326402 270368 326408
rect 270222 5264 270278 5273
rect 270222 5199 270278 5208
rect 270328 4865 270356 326402
rect 270420 5001 270448 335582
rect 270512 328370 270540 335582
rect 270500 328364 270552 328370
rect 270500 328306 270552 328312
rect 270604 326738 270632 340068
rect 270788 340054 270894 340082
rect 270684 339108 270736 339114
rect 270684 339050 270736 339056
rect 270592 326732 270644 326738
rect 270592 326674 270644 326680
rect 270696 326398 270724 339050
rect 270788 326670 270816 340054
rect 271156 339114 271184 340068
rect 271354 340054 271552 340082
rect 271144 339108 271196 339114
rect 271144 339050 271196 339056
rect 271524 335492 271552 340054
rect 271616 335646 271644 340068
rect 271604 335640 271656 335646
rect 271604 335582 271656 335588
rect 271524 335464 271736 335492
rect 271512 328364 271564 328370
rect 271512 328306 271564 328312
rect 270776 326664 270828 326670
rect 270776 326606 270828 326612
rect 271420 326664 271472 326670
rect 271420 326606 271472 326612
rect 270684 326392 270736 326398
rect 270684 326334 270736 326340
rect 271432 11150 271460 326606
rect 271524 11218 271552 328306
rect 271604 326732 271656 326738
rect 271604 326674 271656 326680
rect 271512 11212 271564 11218
rect 271512 11154 271564 11160
rect 271420 11144 271472 11150
rect 271420 11086 271472 11092
rect 271616 9042 271644 326674
rect 271604 9036 271656 9042
rect 271604 8978 271656 8984
rect 271708 8362 271736 335464
rect 271892 326398 271920 340068
rect 271972 336728 272024 336734
rect 271972 336670 272024 336676
rect 271788 326392 271840 326398
rect 271788 326334 271840 326340
rect 271880 326392 271932 326398
rect 271880 326334 271932 326340
rect 271696 8356 271748 8362
rect 271696 8298 271748 8304
rect 271696 6792 271748 6798
rect 271696 6734 271748 6740
rect 270500 5024 270552 5030
rect 270406 4992 270462 5001
rect 270500 4966 270552 4972
rect 270406 4927 270462 4936
rect 270314 4856 270370 4865
rect 270314 4791 270370 4800
rect 270512 480 270540 4966
rect 271708 480 271736 6734
rect 271800 4214 271828 326334
rect 271984 316742 272012 336670
rect 272076 335646 272104 340068
rect 272260 340054 272366 340082
rect 272156 338428 272208 338434
rect 272156 338370 272208 338376
rect 272168 336734 272196 338370
rect 272260 336977 272288 340054
rect 272628 338434 272656 340068
rect 272826 340054 273024 340082
rect 272616 338428 272668 338434
rect 272616 338370 272668 338376
rect 272246 336968 272302 336977
rect 272246 336903 272302 336912
rect 272522 336832 272578 336841
rect 272522 336767 272578 336776
rect 272156 336728 272208 336734
rect 272536 336705 272564 336767
rect 272156 336670 272208 336676
rect 272338 336696 272394 336705
rect 272338 336631 272394 336640
rect 272522 336696 272578 336705
rect 272522 336631 272578 336640
rect 272064 335640 272116 335646
rect 272064 335582 272116 335588
rect 272248 331900 272300 331906
rect 272248 331842 272300 331848
rect 272260 324970 272288 331842
rect 272352 327146 272380 336631
rect 272996 330154 273024 340054
rect 273088 331906 273116 340068
rect 273378 340054 273484 340082
rect 273456 335850 273484 340054
rect 273444 335844 273496 335850
rect 273444 335786 273496 335792
rect 273168 335640 273220 335646
rect 273548 335594 273576 340068
rect 273628 335844 273680 335850
rect 273628 335786 273680 335792
rect 273168 335582 273220 335588
rect 273076 331900 273128 331906
rect 273076 331842 273128 331848
rect 272996 330126 273116 330154
rect 272340 327140 272392 327146
rect 272340 327082 272392 327088
rect 272524 327140 272576 327146
rect 272524 327082 272576 327088
rect 272248 324964 272300 324970
rect 272248 324906 272300 324912
rect 272536 318850 272564 327082
rect 272984 326392 273036 326398
rect 272984 326334 273036 326340
rect 272800 324964 272852 324970
rect 272800 324906 272852 324912
rect 272524 318844 272576 318850
rect 272524 318786 272576 318792
rect 271972 316736 272024 316742
rect 271972 316678 272024 316684
rect 272708 316736 272760 316742
rect 272708 316678 272760 316684
rect 272720 16794 272748 316678
rect 272812 16862 272840 324906
rect 272892 318844 272944 318850
rect 272892 318786 272944 318792
rect 272800 16856 272852 16862
rect 272800 16798 272852 16804
rect 272708 16788 272760 16794
rect 272708 16730 272760 16736
rect 272904 16726 272932 318786
rect 272892 16720 272944 16726
rect 272892 16662 272944 16668
rect 272996 16658 273024 326334
rect 272984 16652 273036 16658
rect 272984 16594 273036 16600
rect 273088 8498 273116 330126
rect 273076 8492 273128 8498
rect 273076 8434 273128 8440
rect 273180 8430 273208 335582
rect 273272 335566 273576 335594
rect 273272 326330 273300 335566
rect 273640 327486 273668 335786
rect 273720 335640 273772 335646
rect 273720 335582 273772 335588
rect 273628 327480 273680 327486
rect 273628 327422 273680 327428
rect 273444 327276 273496 327282
rect 273444 327218 273496 327224
rect 273456 326466 273484 327218
rect 273444 326460 273496 326466
rect 273444 326402 273496 326408
rect 273732 326398 273760 335582
rect 273720 326392 273772 326398
rect 273720 326334 273772 326340
rect 273260 326324 273312 326330
rect 273260 326266 273312 326272
rect 273824 318850 273852 340068
rect 273916 340054 274114 340082
rect 274298 340054 274496 340082
rect 273916 327282 273944 340054
rect 274180 327480 274232 327486
rect 274180 327422 274232 327428
rect 273904 327276 273956 327282
rect 273904 327218 273956 327224
rect 273812 318844 273864 318850
rect 273812 318786 273864 318792
rect 274088 318844 274140 318850
rect 274088 318786 274140 318792
rect 274100 17066 274128 318786
rect 274088 17060 274140 17066
rect 274088 17002 274140 17008
rect 274192 16930 274220 327422
rect 274272 326460 274324 326466
rect 274272 326402 274324 326408
rect 274284 16998 274312 326402
rect 274364 326392 274416 326398
rect 274364 326334 274416 326340
rect 274272 16992 274324 16998
rect 274272 16934 274324 16940
rect 274180 16924 274232 16930
rect 274180 16866 274232 16872
rect 274376 12510 274404 326334
rect 274364 12504 274416 12510
rect 274364 12446 274416 12452
rect 274468 8634 274496 340054
rect 274560 335646 274588 340068
rect 274850 340054 274956 340082
rect 274548 335640 274600 335646
rect 274548 335582 274600 335588
rect 274928 333538 274956 340054
rect 274916 333532 274968 333538
rect 274916 333474 274968 333480
rect 275020 333418 275048 340068
rect 274744 333390 275048 333418
rect 275112 340054 275310 340082
rect 275494 340054 275692 340082
rect 274744 326398 274772 333390
rect 275112 333282 275140 340054
rect 275664 334762 275692 340054
rect 275652 334756 275704 334762
rect 275652 334698 275704 334704
rect 275192 333532 275244 333538
rect 275192 333474 275244 333480
rect 275020 333254 275140 333282
rect 274732 326392 274784 326398
rect 274732 326334 274784 326340
rect 274548 326324 274600 326330
rect 274548 326266 274600 326272
rect 274456 8628 274508 8634
rect 274456 8570 274508 8576
rect 274560 8566 274588 326266
rect 275020 323610 275048 333254
rect 275204 333146 275232 333474
rect 275112 333118 275232 333146
rect 275112 326466 275140 333118
rect 275100 326460 275152 326466
rect 275100 326402 275152 326408
rect 275652 326392 275704 326398
rect 275652 326334 275704 326340
rect 275008 323604 275060 323610
rect 275008 323546 275060 323552
rect 275560 323604 275612 323610
rect 275560 323546 275612 323552
rect 275572 12578 275600 323546
rect 275560 12572 275612 12578
rect 275560 12514 275612 12520
rect 275560 12436 275612 12442
rect 275560 12378 275612 12384
rect 274548 8560 274600 8566
rect 274548 8502 274600 8508
rect 273168 8424 273220 8430
rect 273168 8366 273220 8372
rect 272892 6656 272944 6662
rect 272892 6598 272944 6604
rect 271788 4208 271840 4214
rect 271788 4150 271840 4156
rect 272904 480 272932 6598
rect 275284 6520 275336 6526
rect 275284 6462 275336 6468
rect 274088 4276 274140 4282
rect 274088 4218 274140 4224
rect 273074 4176 273130 4185
rect 273074 4111 273130 4120
rect 273350 4176 273406 4185
rect 273350 4111 273406 4120
rect 273088 3738 273116 4111
rect 273364 3738 273392 4111
rect 273076 3732 273128 3738
rect 273076 3674 273128 3680
rect 273352 3732 273404 3738
rect 273352 3674 273404 3680
rect 274100 480 274128 4218
rect 275192 3392 275244 3398
rect 275192 3334 275244 3340
rect 275204 3233 275232 3334
rect 275190 3224 275246 3233
rect 275190 3159 275246 3168
rect 275296 480 275324 6462
rect 275572 5642 275600 12378
rect 275664 8702 275692 326334
rect 275756 8770 275784 340068
rect 276046 340054 276152 340082
rect 276124 335646 276152 340054
rect 276216 335714 276244 340068
rect 276308 340054 276506 340082
rect 276676 340054 276782 340082
rect 276860 340054 276966 340082
rect 277136 340054 277242 340082
rect 276204 335708 276256 335714
rect 276204 335650 276256 335656
rect 276112 335640 276164 335646
rect 276112 335582 276164 335588
rect 276112 335504 276164 335510
rect 276112 335446 276164 335452
rect 275836 334756 275888 334762
rect 275836 334698 275888 334704
rect 275848 12442 275876 334698
rect 275928 326460 275980 326466
rect 275928 326402 275980 326408
rect 275836 12436 275888 12442
rect 275836 12378 275888 12384
rect 275744 8764 275796 8770
rect 275744 8706 275796 8712
rect 275652 8696 275704 8702
rect 275652 8638 275704 8644
rect 275560 5636 275612 5642
rect 275560 5578 275612 5584
rect 275940 5574 275968 326402
rect 276124 326330 276152 335446
rect 276308 326466 276336 340054
rect 276572 335640 276624 335646
rect 276572 335582 276624 335588
rect 276296 326460 276348 326466
rect 276296 326402 276348 326408
rect 276112 326324 276164 326330
rect 276112 326266 276164 326272
rect 276584 323762 276612 335582
rect 276676 335510 276704 340054
rect 276664 335504 276716 335510
rect 276664 335446 276716 335452
rect 276860 333282 276888 340054
rect 276676 333254 276888 333282
rect 276676 326398 276704 333254
rect 277032 326460 277084 326466
rect 277032 326402 277084 326408
rect 276664 326392 276716 326398
rect 276664 326334 276716 326340
rect 276940 326324 276992 326330
rect 276940 326266 276992 326272
rect 276584 323734 276888 323762
rect 276860 12646 276888 323734
rect 276952 12714 276980 326266
rect 276940 12708 276992 12714
rect 276940 12650 276992 12656
rect 276848 12640 276900 12646
rect 276848 12582 276900 12588
rect 277044 8838 277072 326402
rect 277136 8906 277164 340054
rect 277308 335708 277360 335714
rect 277308 335650 277360 335656
rect 277400 335708 277452 335714
rect 277400 335650 277452 335656
rect 277216 326392 277268 326398
rect 277216 326334 277268 326340
rect 277124 8900 277176 8906
rect 277124 8842 277176 8848
rect 277032 8832 277084 8838
rect 277032 8774 277084 8780
rect 276480 6588 276532 6594
rect 276480 6530 276532 6536
rect 275928 5568 275980 5574
rect 275928 5510 275980 5516
rect 276492 480 276520 6530
rect 277228 5778 277256 326334
rect 277216 5772 277268 5778
rect 277216 5714 277268 5720
rect 277320 5710 277348 335650
rect 277412 326330 277440 335650
rect 277400 326324 277452 326330
rect 277400 326266 277452 326272
rect 277504 323626 277532 340068
rect 277584 335572 277636 335578
rect 277584 335514 277636 335520
rect 277596 328506 277624 335514
rect 277584 328500 277636 328506
rect 277584 328442 277636 328448
rect 277688 326398 277716 340068
rect 277978 340054 278176 340082
rect 277768 335640 277820 335646
rect 277768 335582 277820 335588
rect 277780 326466 277808 335582
rect 278148 335492 278176 340054
rect 278240 335714 278268 340068
rect 278332 340054 278438 340082
rect 278516 340054 278714 340082
rect 278884 340054 278990 340082
rect 279068 340054 279174 340082
rect 279252 340054 279450 340082
rect 278228 335708 278280 335714
rect 278228 335650 278280 335656
rect 278332 335646 278360 340054
rect 278320 335640 278372 335646
rect 278320 335582 278372 335588
rect 278516 335578 278544 340054
rect 278504 335572 278556 335578
rect 278504 335514 278556 335520
rect 278148 335464 278452 335492
rect 277768 326460 277820 326466
rect 277768 326402 277820 326408
rect 277676 326392 277728 326398
rect 277676 326334 277728 326340
rect 278320 326324 278372 326330
rect 278320 326266 278372 326272
rect 277504 323598 277624 323626
rect 277596 321502 277624 323598
rect 277584 321496 277636 321502
rect 277584 321438 277636 321444
rect 278228 321496 278280 321502
rect 278228 321438 278280 321444
rect 278240 17134 278268 321438
rect 278332 17134 278360 326266
rect 278424 17202 278452 335464
rect 278780 334756 278832 334762
rect 278780 334698 278832 334704
rect 278504 328500 278556 328506
rect 278504 328442 278556 328448
rect 278412 17196 278464 17202
rect 278412 17138 278464 17144
rect 278516 17134 278544 328442
rect 278792 326466 278820 334698
rect 278688 326460 278740 326466
rect 278688 326402 278740 326408
rect 278780 326460 278832 326466
rect 278780 326402 278832 326408
rect 278596 326392 278648 326398
rect 278596 326334 278648 326340
rect 278608 17202 278636 326334
rect 278596 17196 278648 17202
rect 278596 17138 278648 17144
rect 278700 17134 278728 326402
rect 278884 326398 278912 340054
rect 278872 326392 278924 326398
rect 278872 326334 278924 326340
rect 279068 326330 279096 340054
rect 279252 334762 279280 340054
rect 279528 336734 279556 340190
rect 281724 340138 281776 340144
rect 282460 340196 282670 340202
rect 282512 340190 282670 340196
rect 299572 340196 299624 340202
rect 282460 340138 282512 340144
rect 299572 340138 299624 340144
rect 300584 340196 300794 340202
rect 300636 340190 300794 340196
rect 305196 340190 305394 340218
rect 317906 340202 318012 340218
rect 317906 340196 318024 340202
rect 317906 340190 317972 340196
rect 300584 340138 300636 340144
rect 279910 340054 280016 340082
rect 279516 336728 279568 336734
rect 279516 336670 279568 336676
rect 279240 334756 279292 334762
rect 279240 334698 279292 334704
rect 279516 327140 279568 327146
rect 279516 327082 279568 327088
rect 279056 326324 279108 326330
rect 279056 326266 279108 326272
rect 279528 323626 279556 327082
rect 279884 326460 279936 326466
rect 279884 326402 279936 326408
rect 279792 326392 279844 326398
rect 279792 326334 279844 326340
rect 279528 323598 279648 323626
rect 279620 321450 279648 323598
rect 279620 321422 279740 321450
rect 278870 63744 278926 63753
rect 278870 63679 278926 63688
rect 278884 63594 278912 63679
rect 278962 63608 279018 63617
rect 278884 63566 278962 63594
rect 278962 63543 279018 63552
rect 278228 17128 278280 17134
rect 278228 17070 278280 17076
rect 278320 17128 278372 17134
rect 278320 17070 278372 17076
rect 278504 17128 278556 17134
rect 278504 17070 278556 17076
rect 278688 17128 278740 17134
rect 278688 17070 278740 17076
rect 278502 16552 278558 16561
rect 278686 16552 278742 16561
rect 278558 16510 278686 16538
rect 278502 16487 278558 16496
rect 278686 16487 278742 16496
rect 278134 16280 278190 16289
rect 278686 16280 278742 16289
rect 278190 16238 278686 16266
rect 278134 16215 278190 16224
rect 278686 16215 278742 16224
rect 278688 13116 278740 13122
rect 278688 13058 278740 13064
rect 278596 12096 278648 12102
rect 278596 12038 278648 12044
rect 278608 5846 278636 12038
rect 278700 5914 278728 13058
rect 279712 12986 279740 321422
rect 279700 12980 279752 12986
rect 279700 12922 279752 12928
rect 279804 12918 279832 326334
rect 279792 12912 279844 12918
rect 279792 12854 279844 12860
rect 279896 9518 279924 326402
rect 279884 9512 279936 9518
rect 279884 9454 279936 9460
rect 278872 6452 278924 6458
rect 278872 6394 278924 6400
rect 278688 5908 278740 5914
rect 278688 5850 278740 5856
rect 278596 5840 278648 5846
rect 278596 5782 278648 5788
rect 277308 5704 277360 5710
rect 277308 5646 277360 5652
rect 277676 4344 277728 4350
rect 277676 4286 277728 4292
rect 277688 480 277716 4286
rect 278884 480 278912 6394
rect 279988 6050 280016 340054
rect 280172 335714 280200 340068
rect 280462 340054 280568 340082
rect 280252 338428 280304 338434
rect 280252 338370 280304 338376
rect 280160 335708 280212 335714
rect 280160 335650 280212 335656
rect 280264 326466 280292 338370
rect 280344 335640 280396 335646
rect 280344 335582 280396 335588
rect 280252 326460 280304 326466
rect 280252 326402 280304 326408
rect 280356 326398 280384 335582
rect 280540 333282 280568 340054
rect 280632 338434 280660 340068
rect 280724 340054 280922 340082
rect 281092 340054 281198 340082
rect 280620 338428 280672 338434
rect 280620 338370 280672 338376
rect 280724 335646 280752 340054
rect 280712 335640 280764 335646
rect 280712 335582 280764 335588
rect 280540 333254 280660 333282
rect 280632 328438 280660 333254
rect 280620 328432 280672 328438
rect 280620 328374 280672 328380
rect 280344 326392 280396 326398
rect 280344 326334 280396 326340
rect 280068 326324 280120 326330
rect 280068 326266 280120 326272
rect 279976 6044 280028 6050
rect 279976 5986 280028 5992
rect 280080 5982 280108 326266
rect 280988 318844 281040 318850
rect 280988 318786 281040 318792
rect 281000 318730 281028 318786
rect 280908 318702 281028 318730
rect 280908 309194 280936 318702
rect 280896 309188 280948 309194
rect 280896 309130 280948 309136
rect 280988 309188 281040 309194
rect 280988 309130 281040 309136
rect 281000 13054 281028 309130
rect 281092 13802 281120 340054
rect 281264 335708 281316 335714
rect 281264 335650 281316 335656
rect 281172 326392 281224 326398
rect 281172 326334 281224 326340
rect 281080 13796 281132 13802
rect 281080 13738 281132 13744
rect 280988 13048 281040 13054
rect 280988 12990 281040 12996
rect 281184 9382 281212 326334
rect 281276 9450 281304 335650
rect 281264 9444 281316 9450
rect 281264 9386 281316 9392
rect 281172 9376 281224 9382
rect 281172 9318 281224 9324
rect 281368 6866 281396 340068
rect 281540 335708 281592 335714
rect 281540 335650 281592 335656
rect 281448 326460 281500 326466
rect 281448 326402 281500 326408
rect 281356 6860 281408 6866
rect 281356 6802 281408 6808
rect 281460 6118 281488 326402
rect 281552 326330 281580 335650
rect 281644 326466 281672 340068
rect 281632 326460 281684 326466
rect 281632 326402 281684 326408
rect 281736 326398 281764 340138
rect 281920 328438 281948 340068
rect 282118 340054 282316 340082
rect 282394 340054 282592 340082
rect 282288 335646 282316 340054
rect 282276 335640 282328 335646
rect 282276 335582 282328 335588
rect 282564 334914 282592 340054
rect 282748 340054 282854 340082
rect 282932 340054 283130 340082
rect 283208 340054 283406 340082
rect 283484 340054 283590 340082
rect 282748 335714 282776 340054
rect 282736 335708 282788 335714
rect 282736 335650 282788 335656
rect 282828 335640 282880 335646
rect 282828 335582 282880 335588
rect 282564 334886 282684 334914
rect 281908 328432 281960 328438
rect 281908 328374 281960 328380
rect 282552 326460 282604 326466
rect 282552 326402 282604 326408
rect 281724 326392 281776 326398
rect 281724 326334 281776 326340
rect 282460 326392 282512 326398
rect 282460 326334 282512 326340
rect 281540 326324 281592 326330
rect 281540 326266 281592 326272
rect 282368 318844 282420 318850
rect 282368 318786 282420 318792
rect 282380 19281 282408 318786
rect 282366 19272 282422 19281
rect 282366 19207 282422 19216
rect 282472 13666 282500 326334
rect 282460 13660 282512 13666
rect 282460 13602 282512 13608
rect 282564 9314 282592 326402
rect 282656 318714 282684 334886
rect 282736 326324 282788 326330
rect 282736 326266 282788 326272
rect 282644 318708 282696 318714
rect 282644 318650 282696 318656
rect 282644 309188 282696 309194
rect 282644 309130 282696 309136
rect 282552 9308 282604 9314
rect 282552 9250 282604 9256
rect 282656 9246 282684 309130
rect 282644 9240 282696 9246
rect 282644 9182 282696 9188
rect 282748 6730 282776 326266
rect 282840 6798 282868 335582
rect 282932 326534 282960 340054
rect 283012 332716 283064 332722
rect 283012 332658 283064 332664
rect 282920 326528 282972 326534
rect 282920 326470 282972 326476
rect 283024 326330 283052 332658
rect 283208 326398 283236 340054
rect 283288 335640 283340 335646
rect 283288 335582 283340 335588
rect 283300 326466 283328 335582
rect 283484 332722 283512 340054
rect 283472 332716 283524 332722
rect 283472 332658 283524 332664
rect 283288 326460 283340 326466
rect 283288 326402 283340 326408
rect 283196 326392 283248 326398
rect 283196 326334 283248 326340
rect 283012 326324 283064 326330
rect 283012 326266 283064 326272
rect 283562 40216 283618 40225
rect 283562 40151 283618 40160
rect 283576 39817 283604 40151
rect 283562 39808 283618 39817
rect 283562 39743 283618 39752
rect 283562 19136 283618 19145
rect 283562 19071 283618 19080
rect 283576 13734 283604 19071
rect 283852 17134 283880 340068
rect 283944 340054 284142 340082
rect 283944 335646 283972 340054
rect 283932 335640 283984 335646
rect 283932 335582 283984 335588
rect 284116 326528 284168 326534
rect 284116 326470 284168 326476
rect 284024 326460 284076 326466
rect 284024 326402 284076 326408
rect 283932 326392 283984 326398
rect 283932 326334 283984 326340
rect 283840 17128 283892 17134
rect 283840 17070 283892 17076
rect 283564 13728 283616 13734
rect 283564 13670 283616 13676
rect 283944 13598 283972 326334
rect 283932 13592 283984 13598
rect 283932 13534 283984 13540
rect 284036 13530 284064 326402
rect 284024 13524 284076 13530
rect 284024 13466 284076 13472
rect 284128 9625 284156 326470
rect 284312 326398 284340 340068
rect 284484 335776 284536 335782
rect 284484 335718 284536 335724
rect 284392 335708 284444 335714
rect 284392 335650 284444 335656
rect 284404 326466 284432 335650
rect 284496 328302 284524 335718
rect 284484 328296 284536 328302
rect 284484 328238 284536 328244
rect 284392 326460 284444 326466
rect 284392 326402 284444 326408
rect 284300 326392 284352 326398
rect 284300 326334 284352 326340
rect 284208 326324 284260 326330
rect 284208 326266 284260 326272
rect 284114 9616 284170 9625
rect 284114 9551 284170 9560
rect 282828 6792 282880 6798
rect 282828 6734 282880 6740
rect 282736 6724 282788 6730
rect 282736 6666 282788 6672
rect 284220 6662 284248 326266
rect 284588 316606 284616 340068
rect 284680 340054 284878 340082
rect 284956 340054 285062 340082
rect 285338 340054 285444 340082
rect 284680 335782 284708 340054
rect 284668 335776 284720 335782
rect 284668 335718 284720 335724
rect 284956 335714 284984 340054
rect 284944 335708 284996 335714
rect 284944 335650 284996 335656
rect 284668 328500 284720 328506
rect 284668 328442 284720 328448
rect 284680 320090 284708 328442
rect 285312 328296 285364 328302
rect 285312 328238 285364 328244
rect 284680 320062 285260 320090
rect 284576 316600 284628 316606
rect 284576 316542 284628 316548
rect 285036 316532 285088 316538
rect 285036 316474 285088 316480
rect 285048 17202 285076 316474
rect 285036 17196 285088 17202
rect 285036 17138 285088 17144
rect 285232 13394 285260 320062
rect 285324 13462 285352 328238
rect 285312 13456 285364 13462
rect 285312 13398 285364 13404
rect 285220 13388 285272 13394
rect 285220 13330 285272 13336
rect 285416 9722 285444 340054
rect 285508 340054 285614 340082
rect 285508 328506 285536 340054
rect 285680 335640 285732 335646
rect 285680 335582 285732 335588
rect 285496 328500 285548 328506
rect 285496 328442 285548 328448
rect 285692 326466 285720 335582
rect 285588 326460 285640 326466
rect 285588 326402 285640 326408
rect 285680 326460 285732 326466
rect 285680 326402 285732 326408
rect 285496 326392 285548 326398
rect 285496 326334 285548 326340
rect 285404 9716 285456 9722
rect 285404 9658 285456 9664
rect 284208 6656 284260 6662
rect 284208 6598 284260 6604
rect 285508 6594 285536 326334
rect 285496 6588 285548 6594
rect 285496 6530 285548 6536
rect 285600 6526 285628 326402
rect 285784 326398 285812 340068
rect 286060 335714 286088 340068
rect 286152 340054 286350 340082
rect 286428 340054 286534 340082
rect 286612 340054 286810 340082
rect 287086 340054 287192 340082
rect 286048 335708 286100 335714
rect 286048 335650 286100 335656
rect 286152 328574 286180 340054
rect 286428 335646 286456 340054
rect 286416 335640 286468 335646
rect 286416 335582 286468 335588
rect 286140 328568 286192 328574
rect 286140 328510 286192 328516
rect 286612 328506 286640 340054
rect 286784 335708 286836 335714
rect 286784 335650 286836 335656
rect 285864 328500 285916 328506
rect 285864 328442 285916 328448
rect 285956 328500 286008 328506
rect 285956 328442 286008 328448
rect 286600 328500 286652 328506
rect 286600 328442 286652 328448
rect 285772 326392 285824 326398
rect 285772 326334 285824 326340
rect 285876 313954 285904 328442
rect 285968 316826 285996 328442
rect 285968 316798 286732 316826
rect 285864 313948 285916 313954
rect 285864 313890 285916 313896
rect 286508 313948 286560 313954
rect 286508 313890 286560 313896
rect 286520 13326 286548 313890
rect 286704 19281 286732 316798
rect 286690 19272 286746 19281
rect 286690 19207 286746 19216
rect 286508 13320 286560 13326
rect 286508 13262 286560 13268
rect 286796 9790 286824 335650
rect 287164 335578 287192 340054
rect 287256 338434 287284 340068
rect 287440 340054 287546 340082
rect 287244 338428 287296 338434
rect 287244 338370 287296 338376
rect 287152 335572 287204 335578
rect 287152 335514 287204 335520
rect 287336 332104 287388 332110
rect 287336 332046 287388 332052
rect 286968 326460 287020 326466
rect 286968 326402 287020 326408
rect 286876 326392 286928 326398
rect 286876 326334 286928 326340
rect 286784 9784 286836 9790
rect 286784 9726 286836 9732
rect 285588 6520 285640 6526
rect 285588 6462 285640 6468
rect 286888 6458 286916 326334
rect 286876 6452 286928 6458
rect 286876 6394 286928 6400
rect 286980 6390 287008 326402
rect 287348 326330 287376 332046
rect 287440 327010 287468 340054
rect 287704 338428 287756 338434
rect 287704 338370 287756 338376
rect 287612 335640 287664 335646
rect 287612 335582 287664 335588
rect 287428 327004 287480 327010
rect 287428 326946 287480 326952
rect 287624 326398 287652 335582
rect 287716 326466 287744 338370
rect 287704 326460 287756 326466
rect 287704 326402 287756 326408
rect 287612 326392 287664 326398
rect 287612 326334 287664 326340
rect 287336 326324 287388 326330
rect 287336 326266 287388 326272
rect 287058 40216 287114 40225
rect 287058 40151 287114 40160
rect 287072 39681 287100 40151
rect 287058 39672 287114 39681
rect 287058 39607 287114 39616
rect 287808 13190 287836 340068
rect 287900 340054 288006 340082
rect 288084 340054 288282 340082
rect 287900 332110 287928 340054
rect 288084 335646 288112 340054
rect 288544 335646 288572 340068
rect 288636 340054 288742 340082
rect 288820 340054 289018 340082
rect 289188 340054 289294 340082
rect 289372 340054 289478 340082
rect 289556 340054 289754 340082
rect 288072 335640 288124 335646
rect 288072 335582 288124 335588
rect 288532 335640 288584 335646
rect 288532 335582 288584 335588
rect 287980 335572 288032 335578
rect 287980 335514 288032 335520
rect 287888 332104 287940 332110
rect 287888 332046 287940 332052
rect 287992 13258 288020 335514
rect 288636 333690 288664 340054
rect 288452 333662 288664 333690
rect 288072 327004 288124 327010
rect 288072 326946 288124 326952
rect 287980 13252 288032 13258
rect 287980 13194 288032 13200
rect 287796 13184 287848 13190
rect 287796 13126 287848 13132
rect 288084 9926 288112 326946
rect 288348 326460 288400 326466
rect 288348 326402 288400 326408
rect 288164 326392 288216 326398
rect 288164 326334 288216 326340
rect 288176 9994 288204 326334
rect 288256 326324 288308 326330
rect 288256 326266 288308 326272
rect 288164 9988 288216 9994
rect 288164 9930 288216 9936
rect 288072 9920 288124 9926
rect 288072 9862 288124 9868
rect 286968 6384 287020 6390
rect 286968 6326 287020 6332
rect 282460 6316 282512 6322
rect 282460 6258 282512 6264
rect 281448 6112 281500 6118
rect 281448 6054 281500 6060
rect 280068 5976 280120 5982
rect 280068 5918 280120 5924
rect 281264 4412 281316 4418
rect 281264 4354 281316 4360
rect 280068 604 280120 610
rect 280068 546 280120 552
rect 280080 480 280108 546
rect 281276 480 281304 4354
rect 282472 480 282500 6258
rect 288268 6254 288296 326266
rect 288360 6322 288388 326402
rect 288452 326330 288480 333662
rect 288624 333600 288676 333606
rect 288624 333542 288676 333548
rect 288636 330546 288664 333542
rect 288624 330540 288676 330546
rect 288624 330482 288676 330488
rect 288820 326466 288848 340054
rect 289084 335640 289136 335646
rect 289084 335582 289136 335588
rect 288900 333532 288952 333538
rect 288900 333474 288952 333480
rect 288808 326460 288860 326466
rect 288808 326402 288860 326408
rect 288912 326398 288940 333474
rect 288900 326392 288952 326398
rect 288900 326334 288952 326340
rect 289096 326346 289124 335582
rect 289188 333606 289216 340054
rect 289176 333600 289228 333606
rect 289176 333542 289228 333548
rect 289372 333418 289400 340054
rect 289556 333538 289584 340054
rect 290016 338434 290044 340068
rect 290004 338428 290056 338434
rect 290004 338370 290056 338376
rect 289912 335708 289964 335714
rect 289912 335650 289964 335656
rect 289820 335640 289872 335646
rect 289820 335582 289872 335588
rect 289544 333532 289596 333538
rect 289544 333474 289596 333480
rect 289188 333390 289400 333418
rect 289188 330664 289216 333390
rect 289188 330636 289492 330664
rect 289360 330540 289412 330546
rect 289360 330482 289412 330488
rect 288440 326324 288492 326330
rect 289096 326318 289308 326346
rect 288440 326266 288492 326272
rect 289280 311982 289308 326318
rect 289268 311976 289320 311982
rect 289268 311918 289320 311924
rect 289176 311840 289228 311846
rect 289176 311782 289228 311788
rect 288438 19136 288494 19145
rect 288438 19071 288494 19080
rect 288452 9858 288480 19071
rect 289188 13122 289216 311782
rect 289372 13705 289400 330482
rect 289464 326754 289492 330636
rect 289464 326726 289676 326754
rect 289544 326460 289596 326466
rect 289544 326402 289596 326408
rect 289452 326392 289504 326398
rect 289452 326334 289504 326340
rect 289358 13696 289414 13705
rect 289358 13631 289414 13640
rect 289176 13116 289228 13122
rect 289176 13058 289228 13064
rect 289464 10130 289492 326334
rect 289452 10124 289504 10130
rect 289452 10066 289504 10072
rect 289556 10062 289584 326402
rect 289544 10056 289596 10062
rect 289544 9998 289596 10004
rect 288440 9852 288492 9858
rect 288440 9794 288492 9800
rect 289648 6769 289676 326726
rect 289832 326330 289860 335582
rect 289924 326534 289952 335650
rect 290096 331084 290148 331090
rect 290096 331026 290148 331032
rect 289912 326528 289964 326534
rect 289912 326470 289964 326476
rect 290108 326466 290136 331026
rect 290096 326460 290148 326466
rect 290096 326402 290148 326408
rect 290200 326398 290228 340068
rect 290384 340054 290490 340082
rect 290568 340054 290674 340082
rect 290752 340054 290950 340082
rect 291226 340054 291332 340082
rect 290280 338428 290332 338434
rect 290280 338370 290332 338376
rect 290292 328438 290320 338370
rect 290384 331090 290412 340054
rect 290568 335646 290596 340054
rect 290752 335714 290780 340054
rect 291304 335782 291332 340054
rect 291396 336666 291424 340068
rect 291384 336660 291436 336666
rect 291384 336602 291436 336608
rect 291292 335776 291344 335782
rect 291292 335718 291344 335724
rect 290740 335708 290792 335714
rect 290740 335650 290792 335656
rect 291568 335708 291620 335714
rect 291568 335650 291620 335656
rect 290556 335640 290608 335646
rect 290556 335582 290608 335588
rect 291476 335640 291528 335646
rect 291476 335582 291528 335588
rect 291292 335572 291344 335578
rect 291292 335514 291344 335520
rect 290372 331084 290424 331090
rect 290372 331026 290424 331032
rect 290280 328432 290332 328438
rect 290280 328374 290332 328380
rect 290648 328432 290700 328438
rect 290648 328374 290700 328380
rect 290188 326392 290240 326398
rect 290188 326334 290240 326340
rect 289728 326324 289780 326330
rect 289728 326266 289780 326272
rect 289820 326324 289872 326330
rect 289820 326266 289872 326272
rect 289634 6760 289690 6769
rect 289634 6695 289690 6704
rect 288348 6316 288400 6322
rect 288348 6258 288400 6264
rect 285956 6248 286008 6254
rect 285956 6190 286008 6196
rect 288256 6248 288308 6254
rect 288256 6190 288308 6196
rect 284760 4548 284812 4554
rect 284760 4490 284812 4496
rect 283656 4480 283708 4486
rect 283656 4422 283708 4428
rect 282828 3596 282880 3602
rect 282828 3538 282880 3544
rect 282840 3233 282868 3538
rect 282826 3224 282882 3233
rect 282826 3159 282882 3168
rect 283668 480 283696 4422
rect 284772 480 284800 4490
rect 285968 480 285996 6190
rect 289740 6186 289768 326266
rect 290660 13569 290688 328374
rect 291304 326534 291332 335514
rect 291108 326528 291160 326534
rect 291108 326470 291160 326476
rect 291292 326528 291344 326534
rect 291292 326470 291344 326476
rect 290924 326460 290976 326466
rect 290924 326402 290976 326408
rect 290832 326324 290884 326330
rect 290832 326266 290884 326272
rect 290646 13560 290702 13569
rect 290646 13495 290702 13504
rect 290844 13433 290872 326266
rect 290830 13424 290886 13433
rect 290830 13359 290886 13368
rect 290936 10198 290964 326402
rect 291016 326392 291068 326398
rect 291016 326334 291068 326340
rect 290924 10192 290976 10198
rect 290924 10134 290976 10140
rect 291028 6633 291056 326334
rect 291014 6624 291070 6633
rect 291014 6559 291070 6568
rect 291120 6497 291148 326470
rect 291488 326466 291516 335582
rect 291476 326460 291528 326466
rect 291476 326402 291528 326408
rect 291580 326398 291608 335650
rect 291568 326392 291620 326398
rect 291568 326334 291620 326340
rect 291672 326330 291700 340068
rect 291856 340054 291962 340082
rect 292040 340054 292146 340082
rect 292224 340054 292422 340082
rect 292592 340054 292698 340082
rect 291752 336660 291804 336666
rect 291752 336602 291804 336608
rect 291764 328438 291792 336602
rect 291856 335646 291884 340054
rect 292040 335714 292068 340054
rect 292028 335708 292080 335714
rect 292028 335650 292080 335656
rect 291844 335640 291896 335646
rect 291844 335582 291896 335588
rect 292224 335578 292252 340054
rect 292304 335776 292356 335782
rect 292304 335718 292356 335724
rect 292212 335572 292264 335578
rect 292212 335514 292264 335520
rect 291752 328432 291804 328438
rect 291752 328374 291804 328380
rect 291936 328432 291988 328438
rect 291936 328374 291988 328380
rect 291660 326324 291712 326330
rect 291660 326266 291712 326272
rect 291948 13297 291976 328374
rect 292212 326460 292264 326466
rect 292212 326402 292264 326408
rect 292120 326392 292172 326398
rect 292120 326334 292172 326340
rect 291934 13288 291990 13297
rect 291934 13223 291990 13232
rect 292132 13161 292160 326334
rect 292118 13152 292174 13161
rect 292118 13087 292174 13096
rect 292224 11014 292252 326402
rect 292212 11008 292264 11014
rect 292212 10950 292264 10956
rect 292316 10266 292344 335718
rect 292488 326528 292540 326534
rect 292488 326470 292540 326476
rect 292396 326324 292448 326330
rect 292396 326266 292448 326272
rect 292304 10260 292356 10266
rect 292304 10202 292356 10208
rect 291106 6488 291162 6497
rect 291106 6423 291162 6432
rect 292408 6361 292436 326266
rect 292394 6352 292450 6361
rect 292394 6287 292450 6296
rect 292500 6225 292528 326470
rect 292592 326262 292620 340054
rect 292764 335572 292816 335578
rect 292764 335514 292816 335520
rect 292776 326534 292804 335514
rect 292764 326528 292816 326534
rect 292764 326470 292816 326476
rect 292868 326330 292896 340068
rect 293158 340054 293356 340082
rect 293040 335708 293092 335714
rect 293040 335650 293092 335656
rect 292948 335640 293000 335646
rect 292948 335582 293000 335588
rect 292960 326466 292988 335582
rect 292948 326460 293000 326466
rect 292948 326402 293000 326408
rect 293052 326398 293080 335650
rect 293040 326392 293092 326398
rect 293040 326334 293092 326340
rect 292856 326324 292908 326330
rect 292856 326266 292908 326272
rect 292580 326256 292632 326262
rect 292580 326198 292632 326204
rect 293328 317490 293356 340054
rect 293420 335578 293448 340068
rect 293512 340054 293618 340082
rect 293696 340054 293894 340082
rect 294064 340054 294170 340082
rect 293512 335646 293540 340054
rect 293696 335714 293724 340054
rect 293684 335708 293736 335714
rect 293684 335650 293736 335656
rect 293500 335640 293552 335646
rect 293500 335582 293552 335588
rect 293408 335572 293460 335578
rect 293408 335514 293460 335520
rect 293960 333328 294012 333334
rect 293960 333270 294012 333276
rect 293776 326528 293828 326534
rect 293776 326470 293828 326476
rect 293592 326460 293644 326466
rect 293592 326402 293644 326408
rect 293500 326392 293552 326398
rect 293500 326334 293552 326340
rect 293316 317484 293368 317490
rect 293316 317426 293368 317432
rect 293408 317484 293460 317490
rect 293408 317426 293460 317432
rect 293420 316010 293448 317426
rect 293328 315982 293448 316010
rect 293328 309194 293356 315982
rect 293316 309188 293368 309194
rect 293316 309130 293368 309136
rect 293408 306400 293460 306406
rect 293408 306342 293460 306348
rect 293420 298178 293448 306342
rect 293316 298172 293368 298178
rect 293316 298114 293368 298120
rect 293408 298172 293460 298178
rect 293408 298114 293460 298120
rect 293328 298058 293356 298114
rect 293236 298030 293356 298058
rect 293236 288454 293264 298030
rect 293224 288448 293276 288454
rect 293130 288416 293186 288425
rect 293316 288448 293368 288454
rect 293224 288390 293276 288396
rect 293314 288416 293316 288425
rect 293368 288416 293370 288425
rect 293130 288351 293186 288360
rect 293314 288351 293370 288360
rect 293144 278798 293172 288351
rect 293132 278792 293184 278798
rect 293132 278734 293184 278740
rect 293316 278792 293368 278798
rect 293316 278734 293368 278740
rect 293328 269113 293356 278734
rect 293130 269104 293186 269113
rect 293130 269039 293186 269048
rect 293314 269104 293370 269113
rect 293314 269039 293370 269048
rect 293144 259486 293172 269039
rect 293132 259480 293184 259486
rect 293132 259422 293184 259428
rect 293316 259480 293368 259486
rect 293316 259422 293368 259428
rect 293328 249801 293356 259422
rect 293130 249792 293186 249801
rect 293130 249727 293186 249736
rect 293314 249792 293370 249801
rect 293314 249727 293370 249736
rect 293144 240174 293172 249727
rect 293132 240168 293184 240174
rect 293132 240110 293184 240116
rect 293316 240168 293368 240174
rect 293316 240110 293368 240116
rect 293328 230489 293356 240110
rect 293130 230480 293186 230489
rect 293130 230415 293186 230424
rect 293314 230480 293370 230489
rect 293314 230415 293370 230424
rect 293144 220862 293172 230415
rect 293132 220856 293184 220862
rect 293130 220824 293132 220833
rect 293316 220856 293368 220862
rect 293184 220824 293186 220833
rect 293130 220759 293186 220768
rect 293314 220824 293316 220833
rect 293368 220824 293370 220833
rect 293314 220759 293370 220768
rect 293144 211177 293172 220759
rect 293130 211168 293186 211177
rect 293130 211103 293132 211112
rect 293184 211103 293186 211112
rect 293314 211168 293370 211177
rect 293314 211103 293316 211112
rect 293132 211074 293184 211080
rect 293368 211103 293370 211112
rect 293316 211074 293368 211080
rect 293144 201521 293172 211074
rect 293130 201512 293186 201521
rect 293130 201447 293132 201456
rect 293184 201447 293186 201456
rect 293314 201512 293370 201521
rect 293314 201447 293316 201456
rect 293132 201418 293184 201424
rect 293368 201447 293370 201456
rect 293316 201418 293368 201424
rect 293144 191865 293172 201418
rect 293130 191856 293186 191865
rect 293130 191791 293132 191800
rect 293184 191791 293186 191800
rect 293314 191856 293370 191865
rect 293314 191791 293316 191800
rect 293132 191762 293184 191768
rect 293368 191791 293370 191800
rect 293316 191762 293368 191768
rect 293144 182209 293172 191762
rect 293130 182200 293186 182209
rect 293130 182135 293132 182144
rect 293184 182135 293186 182144
rect 293314 182200 293370 182209
rect 293314 182135 293316 182144
rect 293132 182106 293184 182112
rect 293368 182135 293370 182144
rect 293316 182106 293368 182112
rect 293144 180810 293172 182106
rect 293132 180804 293184 180810
rect 293132 180746 293184 180752
rect 293316 171148 293368 171154
rect 293316 171090 293368 171096
rect 293328 161430 293356 171090
rect 293316 161424 293368 161430
rect 293316 161366 293368 161372
rect 293316 151836 293368 151842
rect 293316 151778 293368 151784
rect 293328 142118 293356 151778
rect 293316 142112 293368 142118
rect 293316 142054 293368 142060
rect 293316 132524 293368 132530
rect 293316 132466 293368 132472
rect 293328 103494 293356 132466
rect 293316 103488 293368 103494
rect 293316 103430 293368 103436
rect 293316 93900 293368 93906
rect 293316 93842 293368 93848
rect 293328 84182 293356 93842
rect 293316 84176 293368 84182
rect 293316 84118 293368 84124
rect 293316 74588 293368 74594
rect 293316 74530 293368 74536
rect 293328 64870 293356 74530
rect 293316 64864 293368 64870
rect 293316 64806 293368 64812
rect 293408 46980 293460 46986
rect 293408 46922 293460 46928
rect 293420 17882 293448 46922
rect 293408 17876 293460 17882
rect 293408 17818 293460 17824
rect 293512 17746 293540 326334
rect 293604 17814 293632 326402
rect 293684 326324 293736 326330
rect 293684 326266 293736 326272
rect 293696 17950 293724 326266
rect 293684 17944 293736 17950
rect 293684 17886 293736 17892
rect 293592 17808 293644 17814
rect 293592 17750 293644 17756
rect 293500 17740 293552 17746
rect 293500 17682 293552 17688
rect 292578 17096 292634 17105
rect 292578 17031 292634 17040
rect 292592 16833 292620 17031
rect 292578 16824 292634 16833
rect 292578 16759 292634 16768
rect 293788 10878 293816 326470
rect 293868 326256 293920 326262
rect 293868 326198 293920 326204
rect 293880 10946 293908 326198
rect 293972 317490 294000 333270
rect 294064 326466 294092 340054
rect 294236 333192 294288 333198
rect 294236 333134 294288 333140
rect 294052 326460 294104 326466
rect 294052 326402 294104 326408
rect 294248 326398 294276 333134
rect 294236 326392 294288 326398
rect 294236 326334 294288 326340
rect 294340 326346 294368 340068
rect 294432 340054 294630 340082
rect 294906 340054 295012 340082
rect 294432 333198 294460 340054
rect 294420 333192 294472 333198
rect 294420 333134 294472 333140
rect 294984 331242 295012 340054
rect 295076 333334 295104 340068
rect 295064 333328 295116 333334
rect 295064 333270 295116 333276
rect 294984 331214 295196 331242
rect 295064 326392 295116 326398
rect 294340 326318 295012 326346
rect 295064 326334 295116 326340
rect 293960 317484 294012 317490
rect 293960 317426 294012 317432
rect 294788 317484 294840 317490
rect 294788 317426 294840 317432
rect 294800 211313 294828 317426
rect 294786 211304 294842 211313
rect 294786 211239 294842 211248
rect 294786 211168 294842 211177
rect 294604 211132 294656 211138
rect 294786 211103 294788 211112
rect 294604 211074 294656 211080
rect 294840 211103 294842 211112
rect 294788 211074 294840 211080
rect 294616 201521 294644 211074
rect 294602 201512 294658 201521
rect 294602 201447 294658 201456
rect 294786 201512 294842 201521
rect 294786 201447 294842 201456
rect 294800 192001 294828 201447
rect 294786 191992 294842 192001
rect 294786 191927 294842 191936
rect 294786 191856 294842 191865
rect 294604 191820 294656 191826
rect 294786 191791 294788 191800
rect 294604 191762 294656 191768
rect 294840 191791 294842 191800
rect 294788 191762 294840 191768
rect 294616 182209 294644 191762
rect 294602 182200 294658 182209
rect 294602 182135 294658 182144
rect 294786 182200 294842 182209
rect 294786 182135 294842 182144
rect 294800 171290 294828 182135
rect 294788 171284 294840 171290
rect 294788 171226 294840 171232
rect 294788 171148 294840 171154
rect 294788 171090 294840 171096
rect 294800 151978 294828 171090
rect 294788 151972 294840 151978
rect 294788 151914 294840 151920
rect 294788 151836 294840 151842
rect 294788 151778 294840 151784
rect 294800 151722 294828 151778
rect 294708 151694 294828 151722
rect 294708 142186 294736 151694
rect 294696 142180 294748 142186
rect 294696 142122 294748 142128
rect 294788 142180 294840 142186
rect 294788 142122 294840 142128
rect 294800 132818 294828 142122
rect 294800 132790 294920 132818
rect 294892 132530 294920 132790
rect 294788 132524 294840 132530
rect 294788 132466 294840 132472
rect 294880 132524 294932 132530
rect 294880 132466 294932 132472
rect 294800 132410 294828 132466
rect 294708 132382 294828 132410
rect 294708 122874 294736 132382
rect 294696 122868 294748 122874
rect 294696 122810 294748 122816
rect 294788 122868 294840 122874
rect 294788 122810 294840 122816
rect 294800 113150 294828 122810
rect 294788 113144 294840 113150
rect 294788 113086 294840 113092
rect 294788 103556 294840 103562
rect 294788 103498 294840 103504
rect 294800 95334 294828 103498
rect 294788 95328 294840 95334
rect 294788 95270 294840 95276
rect 294696 95192 294748 95198
rect 294696 95134 294748 95140
rect 294708 85610 294736 95134
rect 294696 85604 294748 85610
rect 294696 85546 294748 85552
rect 294788 85604 294840 85610
rect 294788 85546 294840 85552
rect 294800 84182 294828 85546
rect 294788 84176 294840 84182
rect 294788 84118 294840 84124
rect 294788 74588 294840 74594
rect 294788 74530 294840 74536
rect 294800 64870 294828 74530
rect 294788 64864 294840 64870
rect 294788 64806 294840 64812
rect 294880 46980 294932 46986
rect 294880 46922 294932 46928
rect 294892 18562 294920 46922
rect 294880 18556 294932 18562
rect 294880 18498 294932 18504
rect 294984 17678 295012 326318
rect 294972 17672 295024 17678
rect 294972 17614 295024 17620
rect 295076 17610 295104 326334
rect 295064 17604 295116 17610
rect 295064 17546 295116 17552
rect 293868 10940 293920 10946
rect 293868 10882 293920 10888
rect 293776 10872 293828 10878
rect 293776 10814 293828 10820
rect 295168 10742 295196 331214
rect 295248 326460 295300 326466
rect 295248 326402 295300 326408
rect 295260 10810 295288 326402
rect 295352 326398 295380 340068
rect 295444 340054 295642 340082
rect 295720 340054 295826 340082
rect 295904 340054 296102 340082
rect 296378 340054 296484 340082
rect 295444 328778 295472 340054
rect 295616 330880 295668 330886
rect 295616 330822 295668 330828
rect 295432 328772 295484 328778
rect 295432 328714 295484 328720
rect 295628 327078 295656 330822
rect 295616 327072 295668 327078
rect 295616 327014 295668 327020
rect 295340 326392 295392 326398
rect 295340 326334 295392 326340
rect 295720 326346 295748 340054
rect 295904 326466 295932 340054
rect 296352 328772 296404 328778
rect 296352 328714 296404 328720
rect 295892 326460 295944 326466
rect 295892 326402 295944 326408
rect 295720 326318 296300 326346
rect 296076 322244 296128 322250
rect 296076 322186 296128 322192
rect 296088 211313 296116 322186
rect 296074 211304 296130 211313
rect 296074 211239 296130 211248
rect 296074 211168 296130 211177
rect 295892 211132 295944 211138
rect 296074 211103 296076 211112
rect 295892 211074 295944 211080
rect 296128 211103 296130 211112
rect 296076 211074 296128 211080
rect 295904 201521 295932 211074
rect 295890 201512 295946 201521
rect 295890 201447 295946 201456
rect 296074 201512 296130 201521
rect 296074 201447 296130 201456
rect 296088 192001 296116 201447
rect 296074 191992 296130 192001
rect 296074 191927 296130 191936
rect 296074 191856 296130 191865
rect 295892 191820 295944 191826
rect 296074 191791 296076 191800
rect 295892 191762 295944 191768
rect 296128 191791 296130 191800
rect 296076 191762 296128 191768
rect 295904 182209 295932 191762
rect 295890 182200 295946 182209
rect 295890 182135 295946 182144
rect 296074 182200 296130 182209
rect 296074 182135 296130 182144
rect 296088 171290 296116 182135
rect 296076 171284 296128 171290
rect 296076 171226 296128 171232
rect 296076 171148 296128 171154
rect 296076 171090 296128 171096
rect 296088 151978 296116 171090
rect 296076 151972 296128 151978
rect 296076 151914 296128 151920
rect 296076 151836 296128 151842
rect 296076 151778 296128 151784
rect 296088 150414 296116 151778
rect 296076 150408 296128 150414
rect 296076 150350 296128 150356
rect 296168 140820 296220 140826
rect 296168 140762 296220 140768
rect 296180 134586 296208 140762
rect 296088 134558 296208 134586
rect 296088 113098 296116 134558
rect 295996 113070 296116 113098
rect 295996 103562 296024 113070
rect 295984 103556 296036 103562
rect 295984 103498 296036 103504
rect 296076 103556 296128 103562
rect 296076 103498 296128 103504
rect 296088 103442 296116 103498
rect 295996 103414 296116 103442
rect 295996 93906 296024 103414
rect 295984 93900 296036 93906
rect 295984 93842 296036 93848
rect 296076 93900 296128 93906
rect 296076 93842 296128 93848
rect 296088 84130 296116 93842
rect 295996 84102 296116 84130
rect 295996 74594 296024 84102
rect 295984 74588 296036 74594
rect 295984 74530 296036 74536
rect 296076 74588 296128 74594
rect 296076 74530 296128 74536
rect 296088 64818 296116 74530
rect 296088 64790 296208 64818
rect 296180 60042 296208 64790
rect 296168 60036 296220 60042
rect 296168 59978 296220 59984
rect 296168 46980 296220 46986
rect 296168 46922 296220 46928
rect 296180 13938 296208 46922
rect 296168 13932 296220 13938
rect 296168 13874 296220 13880
rect 296272 13870 296300 326318
rect 296260 13864 296312 13870
rect 296260 13806 296312 13812
rect 295248 10804 295300 10810
rect 295248 10746 295300 10752
rect 295156 10736 295208 10742
rect 295156 10678 295208 10684
rect 296364 10674 296392 328714
rect 296352 10668 296404 10674
rect 296352 10610 296404 10616
rect 296456 10606 296484 340054
rect 296548 330886 296576 340068
rect 296824 335714 296852 340068
rect 296916 340054 297114 340082
rect 297192 340054 297298 340082
rect 297376 340054 297574 340082
rect 296812 335708 296864 335714
rect 296812 335650 296864 335656
rect 296916 335594 296944 340054
rect 297192 335696 297220 340054
rect 296732 335566 296944 335594
rect 297008 335668 297220 335696
rect 296536 330880 296588 330886
rect 296536 330822 296588 330828
rect 296536 326460 296588 326466
rect 296536 326402 296588 326408
rect 296444 10600 296496 10606
rect 296444 10542 296496 10548
rect 293132 7948 293184 7954
rect 293132 7890 293184 7896
rect 292486 6216 292542 6225
rect 289544 6180 289596 6186
rect 289544 6122 289596 6128
rect 289728 6180 289780 6186
rect 292486 6151 292542 6160
rect 289728 6122 289780 6128
rect 287152 4684 287204 4690
rect 287152 4626 287204 4632
rect 287164 480 287192 4626
rect 288348 4616 288400 4622
rect 288348 4558 288400 4564
rect 288360 480 288388 4558
rect 289556 480 289584 6122
rect 291936 5500 291988 5506
rect 291936 5442 291988 5448
rect 290740 4752 290792 4758
rect 290740 4694 290792 4700
rect 290752 480 290780 4694
rect 291948 480 291976 5442
rect 292316 4282 292528 4298
rect 292304 4276 292528 4282
rect 292356 4270 292528 4276
rect 292304 4218 292356 4224
rect 292394 4176 292450 4185
rect 292394 4111 292450 4120
rect 292408 3738 292436 4111
rect 292500 3738 292528 4270
rect 292670 4176 292726 4185
rect 292670 4111 292726 4120
rect 292684 3738 292712 4111
rect 292396 3732 292448 3738
rect 292396 3674 292448 3680
rect 292488 3732 292540 3738
rect 292488 3674 292540 3680
rect 292672 3732 292724 3738
rect 292672 3674 292724 3680
rect 293144 480 293172 7890
rect 296548 7138 296576 326402
rect 296732 326398 296760 335566
rect 297008 335458 297036 335668
rect 297376 335594 297404 340054
rect 297456 335708 297508 335714
rect 297456 335650 297508 335656
rect 296916 335430 297036 335458
rect 297192 335566 297404 335594
rect 296628 326392 296680 326398
rect 296628 326334 296680 326340
rect 296720 326392 296772 326398
rect 296720 326334 296772 326340
rect 296640 89078 296668 326334
rect 296916 325582 296944 335430
rect 296996 335368 297048 335374
rect 296996 335310 297048 335316
rect 297008 326380 297036 335310
rect 297192 326602 297220 335566
rect 297468 335458 297496 335650
rect 297376 335430 297496 335458
rect 297180 326596 297232 326602
rect 297180 326538 297232 326544
rect 297376 326534 297404 335430
rect 297364 326528 297416 326534
rect 297364 326470 297416 326476
rect 297732 326392 297784 326398
rect 297008 326352 297680 326380
rect 296904 325576 296956 325582
rect 296904 325518 296956 325524
rect 297548 325576 297600 325582
rect 297548 325518 297600 325524
rect 297560 106962 297588 325518
rect 297548 106956 297600 106962
rect 297548 106898 297600 106904
rect 297456 100768 297508 100774
rect 297456 100710 297508 100716
rect 297468 96694 297496 100710
rect 297456 96688 297508 96694
rect 297456 96630 297508 96636
rect 297548 96552 297600 96558
rect 297548 96494 297600 96500
rect 296628 89072 296680 89078
rect 296628 89014 296680 89020
rect 296628 86896 296680 86902
rect 296628 86838 296680 86844
rect 296536 7132 296588 7138
rect 296536 7074 296588 7080
rect 296640 7070 296668 86838
rect 297560 23390 297588 96494
rect 297652 23458 297680 326352
rect 297732 326334 297784 326340
rect 297640 23452 297692 23458
rect 297640 23394 297692 23400
rect 297548 23384 297600 23390
rect 297548 23326 297600 23332
rect 297362 16280 297418 16289
rect 297362 16215 297418 16224
rect 297376 15609 297404 16215
rect 297362 15600 297418 15609
rect 297362 15535 297418 15544
rect 297744 10538 297772 326334
rect 297732 10532 297784 10538
rect 297732 10474 297784 10480
rect 297836 10470 297864 340068
rect 297928 340054 298034 340082
rect 298310 340054 298416 340082
rect 298586 340054 298692 340082
rect 297928 335374 297956 340054
rect 297916 335368 297968 335374
rect 297916 335310 297968 335316
rect 298100 332784 298152 332790
rect 298100 332726 298152 332732
rect 297916 326596 297968 326602
rect 297916 326538 297968 326544
rect 297824 10464 297876 10470
rect 297824 10406 297876 10412
rect 296720 7880 296772 7886
rect 296720 7822 296772 7828
rect 296628 7064 296680 7070
rect 296628 7006 296680 7012
rect 294328 5432 294380 5438
rect 294328 5374 294380 5380
rect 294340 480 294368 5374
rect 295524 5364 295576 5370
rect 295524 5306 295576 5312
rect 295536 480 295564 5306
rect 296732 480 296760 7822
rect 297928 7274 297956 326538
rect 298008 326528 298060 326534
rect 298008 326470 298060 326476
rect 297916 7268 297968 7274
rect 297916 7210 297968 7216
rect 298020 7206 298048 326470
rect 298112 323474 298140 332726
rect 298192 331424 298244 331430
rect 298192 331366 298244 331372
rect 298204 326466 298232 331366
rect 298192 326460 298244 326466
rect 298192 326402 298244 326408
rect 298388 326398 298416 340054
rect 298468 335640 298520 335646
rect 298468 335582 298520 335588
rect 298376 326392 298428 326398
rect 298376 326334 298428 326340
rect 298480 323610 298508 335582
rect 298664 331650 298692 340054
rect 298756 332790 298784 340068
rect 298848 340054 299046 340082
rect 299124 340054 299322 340082
rect 298744 332784 298796 332790
rect 298744 332726 298796 332732
rect 298664 331622 298784 331650
rect 298756 331158 298784 331622
rect 298848 331430 298876 340054
rect 299124 335646 299152 340054
rect 299112 335640 299164 335646
rect 299112 335582 299164 335588
rect 298836 331424 298888 331430
rect 298836 331366 298888 331372
rect 298744 331152 298796 331158
rect 298744 331094 298796 331100
rect 299204 331152 299256 331158
rect 299204 331094 299256 331100
rect 298468 323604 298520 323610
rect 298468 323546 298520 323552
rect 299112 323604 299164 323610
rect 299112 323546 299164 323552
rect 298100 323468 298152 323474
rect 298100 323410 298152 323416
rect 299020 323468 299072 323474
rect 299020 323410 299072 323416
rect 299032 256698 299060 323410
rect 299020 256692 299072 256698
rect 299020 256634 299072 256640
rect 299020 247104 299072 247110
rect 299020 247046 299072 247052
rect 299032 237386 299060 247046
rect 299020 237380 299072 237386
rect 299020 237322 299072 237328
rect 299020 227792 299072 227798
rect 299020 227734 299072 227740
rect 299032 227662 299060 227734
rect 299020 227656 299072 227662
rect 299020 227598 299072 227604
rect 299020 218068 299072 218074
rect 299020 218010 299072 218016
rect 299032 208554 299060 218010
rect 299020 208548 299072 208554
rect 299020 208490 299072 208496
rect 299020 208412 299072 208418
rect 299020 208354 299072 208360
rect 299032 198694 299060 208354
rect 299020 198688 299072 198694
rect 299020 198630 299072 198636
rect 299020 189100 299072 189106
rect 299020 189042 299072 189048
rect 299032 188986 299060 189042
rect 298940 188958 299060 188986
rect 298940 179450 298968 188958
rect 298928 179444 298980 179450
rect 298928 179386 298980 179392
rect 299020 179444 299072 179450
rect 299020 179386 299072 179392
rect 299032 169726 299060 179386
rect 299020 169720 299072 169726
rect 299020 169662 299072 169668
rect 299020 160132 299072 160138
rect 299020 160074 299072 160080
rect 299032 140758 299060 160074
rect 299020 140752 299072 140758
rect 299020 140694 299072 140700
rect 299020 129872 299072 129878
rect 299020 129814 299072 129820
rect 299032 129742 299060 129814
rect 299020 129736 299072 129742
rect 299020 129678 299072 129684
rect 299020 120216 299072 120222
rect 299020 120158 299072 120164
rect 299032 120086 299060 120158
rect 299020 120080 299072 120086
rect 299020 120022 299072 120028
rect 298928 102196 298980 102202
rect 298928 102138 298980 102144
rect 298940 93838 298968 102138
rect 298928 93832 298980 93838
rect 298928 93774 298980 93780
rect 299020 93764 299072 93770
rect 299020 93706 299072 93712
rect 299032 55214 299060 93706
rect 299020 55208 299072 55214
rect 299020 55150 299072 55156
rect 299020 45620 299072 45626
rect 299020 45562 299072 45568
rect 299032 35902 299060 45562
rect 299020 35896 299072 35902
rect 299020 35838 299072 35844
rect 299020 26308 299072 26314
rect 299020 26250 299072 26256
rect 299032 14142 299060 26250
rect 299020 14136 299072 14142
rect 299020 14078 299072 14084
rect 299124 10334 299152 323546
rect 299216 10402 299244 331094
rect 299388 326460 299440 326466
rect 299388 326402 299440 326408
rect 299296 326392 299348 326398
rect 299296 326334 299348 326340
rect 299204 10396 299256 10402
rect 299204 10338 299256 10344
rect 299112 10328 299164 10334
rect 299112 10270 299164 10276
rect 299308 7342 299336 326334
rect 299400 7410 299428 326402
rect 299492 326194 299520 340068
rect 299480 326188 299532 326194
rect 299480 326130 299532 326136
rect 299584 326126 299612 340138
rect 299664 335844 299716 335850
rect 299664 335786 299716 335792
rect 299676 326262 299704 335786
rect 299768 333282 299796 340068
rect 299860 340054 300058 340082
rect 300136 340054 300242 340082
rect 300518 340054 300716 340082
rect 299860 335850 299888 340054
rect 299848 335844 299900 335850
rect 299848 335786 299900 335792
rect 299768 333254 299980 333282
rect 299848 328568 299900 328574
rect 299848 328510 299900 328516
rect 299664 326256 299716 326262
rect 299664 326198 299716 326204
rect 299572 326120 299624 326126
rect 299572 326062 299624 326068
rect 299860 320906 299888 328510
rect 299952 326346 299980 333254
rect 300136 328574 300164 340054
rect 300688 333690 300716 340054
rect 300872 340054 300978 340082
rect 300688 333662 300808 333690
rect 300124 328568 300176 328574
rect 300124 328510 300176 328516
rect 299952 326318 300716 326346
rect 300492 326256 300544 326262
rect 300492 326198 300544 326204
rect 300400 326188 300452 326194
rect 300400 326130 300452 326136
rect 299860 320878 300256 320906
rect 300228 316044 300256 320878
rect 300228 316016 300348 316044
rect 300320 247042 300348 316016
rect 300308 247036 300360 247042
rect 300308 246978 300360 246984
rect 300308 237448 300360 237454
rect 300308 237390 300360 237396
rect 300320 227730 300348 237390
rect 300308 227724 300360 227730
rect 300308 227666 300360 227672
rect 300308 218068 300360 218074
rect 300308 218010 300360 218016
rect 300320 208350 300348 218010
rect 300308 208344 300360 208350
rect 300308 208286 300360 208292
rect 300308 198756 300360 198762
rect 300308 198698 300360 198704
rect 300320 189038 300348 198698
rect 300308 189032 300360 189038
rect 300308 188974 300360 188980
rect 300308 179444 300360 179450
rect 300308 179386 300360 179392
rect 300320 169726 300348 179386
rect 300308 169720 300360 169726
rect 300308 169662 300360 169668
rect 300308 160132 300360 160138
rect 300308 160074 300360 160080
rect 300320 140758 300348 160074
rect 300308 140752 300360 140758
rect 300308 140694 300360 140700
rect 300308 130756 300360 130762
rect 300308 130698 300360 130704
rect 300320 120086 300348 130698
rect 300308 120080 300360 120086
rect 300308 120022 300360 120028
rect 300216 102196 300268 102202
rect 300216 102138 300268 102144
rect 300228 93838 300256 102138
rect 300216 93832 300268 93838
rect 300216 93774 300268 93780
rect 300308 93764 300360 93770
rect 300308 93706 300360 93712
rect 300320 55214 300348 93706
rect 300308 55208 300360 55214
rect 300308 55150 300360 55156
rect 300308 45620 300360 45626
rect 300308 45562 300360 45568
rect 300320 35902 300348 45562
rect 300308 35896 300360 35902
rect 300308 35838 300360 35844
rect 300308 26308 300360 26314
rect 300308 26250 300360 26256
rect 300320 14278 300348 26250
rect 300308 14272 300360 14278
rect 300308 14214 300360 14220
rect 300412 14210 300440 326130
rect 300400 14204 300452 14210
rect 300400 14146 300452 14152
rect 300504 10849 300532 326198
rect 300584 326120 300636 326126
rect 300584 326062 300636 326068
rect 300490 10840 300546 10849
rect 300490 10775 300546 10784
rect 300596 10713 300624 326062
rect 300582 10704 300638 10713
rect 300582 10639 300638 10648
rect 300308 7812 300360 7818
rect 300308 7754 300360 7760
rect 299388 7404 299440 7410
rect 299388 7346 299440 7352
rect 299296 7336 299348 7342
rect 299296 7278 299348 7284
rect 298008 7200 298060 7206
rect 298008 7142 298060 7148
rect 297916 5296 297968 5302
rect 297916 5238 297968 5244
rect 297928 480 297956 5238
rect 299112 5228 299164 5234
rect 299112 5170 299164 5176
rect 299124 480 299152 5170
rect 300320 480 300348 7754
rect 300688 7478 300716 326318
rect 300780 7546 300808 333662
rect 300872 326262 300900 340054
rect 301240 331362 301268 340068
rect 301332 340054 301530 340082
rect 301608 340054 301714 340082
rect 301990 340054 302096 340082
rect 301228 331356 301280 331362
rect 301228 331298 301280 331304
rect 301332 331242 301360 340054
rect 301056 331214 301360 331242
rect 301056 331140 301084 331214
rect 301056 331112 301176 331140
rect 301044 328568 301096 328574
rect 301044 328510 301096 328516
rect 300860 326256 300912 326262
rect 300860 326198 300912 326204
rect 301056 316062 301084 328510
rect 301148 326346 301176 331112
rect 301228 331084 301280 331090
rect 301228 331026 301280 331032
rect 301240 326466 301268 331026
rect 301608 328574 301636 340054
rect 301596 328568 301648 328574
rect 301596 328510 301648 328516
rect 301228 326460 301280 326466
rect 301228 326402 301280 326408
rect 301148 326318 302004 326346
rect 301872 326256 301924 326262
rect 301872 326198 301924 326204
rect 301044 316056 301096 316062
rect 301044 315998 301096 316004
rect 301780 316056 301832 316062
rect 301780 315998 301832 316004
rect 301792 247042 301820 315998
rect 301780 247036 301832 247042
rect 301780 246978 301832 246984
rect 301780 237448 301832 237454
rect 301780 237390 301832 237396
rect 301792 235958 301820 237390
rect 301780 235952 301832 235958
rect 301780 235894 301832 235900
rect 301780 226364 301832 226370
rect 301780 226306 301832 226312
rect 301792 218362 301820 226306
rect 301608 218334 301820 218362
rect 301608 218113 301636 218334
rect 301594 218104 301650 218113
rect 301594 218039 301650 218048
rect 301778 218104 301834 218113
rect 301778 218039 301834 218048
rect 301792 216646 301820 218039
rect 301780 216640 301832 216646
rect 301780 216582 301832 216588
rect 301596 207052 301648 207058
rect 301596 206994 301648 207000
rect 301608 198801 301636 206994
rect 301594 198792 301650 198801
rect 301594 198727 301650 198736
rect 301778 198792 301834 198801
rect 301778 198727 301834 198736
rect 301792 197334 301820 198727
rect 301780 197328 301832 197334
rect 301780 197270 301832 197276
rect 301780 187740 301832 187746
rect 301780 187682 301832 187688
rect 301792 179654 301820 187682
rect 301780 179648 301832 179654
rect 301780 179590 301832 179596
rect 301780 179512 301832 179518
rect 301780 179454 301832 179460
rect 301792 178022 301820 179454
rect 301780 178016 301832 178022
rect 301780 177958 301832 177964
rect 301780 168428 301832 168434
rect 301780 168370 301832 168376
rect 301792 160138 301820 168370
rect 301884 160410 301912 326198
rect 301872 160404 301924 160410
rect 301872 160346 301924 160352
rect 301780 160132 301832 160138
rect 301780 160074 301832 160080
rect 301872 160132 301924 160138
rect 301872 160074 301924 160080
rect 301780 159996 301832 160002
rect 301780 159938 301832 159944
rect 301792 150278 301820 159938
rect 301780 150272 301832 150278
rect 301780 150214 301832 150220
rect 301504 147688 301556 147694
rect 301504 147630 301556 147636
rect 301516 140758 301544 147630
rect 301884 141098 301912 160074
rect 301976 141273 302004 326318
rect 301962 141264 302018 141273
rect 301962 141199 302018 141208
rect 301872 141092 301924 141098
rect 301872 141034 301924 141040
rect 301962 140856 302018 140865
rect 301962 140791 302018 140800
rect 301504 140752 301556 140758
rect 301504 140694 301556 140700
rect 301780 140752 301832 140758
rect 301780 140694 301832 140700
rect 301792 134570 301820 140694
rect 301872 140684 301924 140690
rect 301872 140626 301924 140632
rect 301780 134564 301832 134570
rect 301780 134506 301832 134512
rect 301780 121508 301832 121514
rect 301780 121450 301832 121456
rect 301792 120086 301820 121450
rect 301780 120080 301832 120086
rect 301780 120022 301832 120028
rect 301688 102196 301740 102202
rect 301688 102138 301740 102144
rect 301700 93838 301728 102138
rect 301688 93832 301740 93838
rect 301688 93774 301740 93780
rect 301780 93764 301832 93770
rect 301780 93706 301832 93712
rect 301792 55214 301820 93706
rect 301780 55208 301832 55214
rect 301780 55150 301832 55156
rect 301780 45620 301832 45626
rect 301780 45562 301832 45568
rect 301792 35902 301820 45562
rect 301780 35896 301832 35902
rect 301780 35838 301832 35844
rect 301780 26308 301832 26314
rect 301780 26250 301832 26256
rect 301792 18290 301820 26250
rect 301780 18284 301832 18290
rect 301780 18226 301832 18232
rect 301884 18222 301912 140626
rect 301872 18216 301924 18222
rect 301872 18158 301924 18164
rect 301976 17270 302004 140791
rect 302068 17338 302096 340054
rect 302252 326466 302280 340068
rect 302344 340054 302450 340082
rect 302344 330614 302372 340054
rect 302608 335640 302660 335646
rect 302608 335582 302660 335588
rect 302332 330608 302384 330614
rect 302332 330550 302384 330556
rect 302148 326460 302200 326466
rect 302148 326402 302200 326408
rect 302240 326460 302292 326466
rect 302240 326402 302292 326408
rect 302056 17332 302108 17338
rect 302056 17274 302108 17280
rect 302160 17270 302188 326402
rect 302620 321502 302648 335582
rect 302712 326398 302740 340068
rect 302988 339114 303016 340068
rect 303186 340054 303292 340082
rect 302976 339108 303028 339114
rect 302976 339050 303028 339056
rect 303160 330608 303212 330614
rect 303160 330550 303212 330556
rect 302700 326392 302752 326398
rect 302700 326334 302752 326340
rect 302608 321496 302660 321502
rect 302608 321438 302660 321444
rect 303068 321496 303120 321502
rect 303068 321438 303120 321444
rect 303080 17542 303108 321438
rect 303068 17536 303120 17542
rect 303068 17478 303120 17484
rect 301964 17264 302016 17270
rect 301964 17206 302016 17212
rect 302148 17264 302200 17270
rect 302148 17206 302200 17212
rect 300858 17096 300914 17105
rect 300858 17031 300914 17040
rect 300872 16969 300900 17031
rect 300858 16960 300914 16969
rect 300858 16895 300914 16904
rect 301964 15224 302016 15230
rect 301964 15166 302016 15172
rect 302148 15224 302200 15230
rect 302148 15166 302200 15172
rect 301976 10577 302004 15166
rect 302056 15156 302108 15162
rect 302056 15098 302108 15104
rect 301962 10568 302018 10577
rect 301962 10503 302018 10512
rect 302068 8226 302096 15098
rect 302160 8294 302188 15166
rect 303172 15162 303200 330550
rect 303160 15156 303212 15162
rect 303160 15098 303212 15104
rect 303264 15094 303292 340054
rect 303344 339108 303396 339114
rect 303344 339050 303396 339056
rect 303252 15088 303304 15094
rect 303252 15030 303304 15036
rect 303356 10305 303384 339050
rect 303448 335646 303476 340068
rect 303632 340054 303738 340082
rect 303436 335640 303488 335646
rect 303436 335582 303488 335588
rect 303436 326460 303488 326466
rect 303436 326402 303488 326408
rect 303448 10441 303476 326402
rect 303528 326392 303580 326398
rect 303528 326334 303580 326340
rect 303434 10432 303490 10441
rect 303434 10367 303490 10376
rect 303342 10296 303398 10305
rect 303342 10231 303398 10240
rect 302148 8288 302200 8294
rect 302148 8230 302200 8236
rect 302056 8220 302108 8226
rect 302056 8162 302108 8168
rect 303540 8158 303568 326334
rect 303632 326330 303660 340054
rect 303804 335776 303856 335782
rect 303804 335718 303856 335724
rect 303816 326398 303844 335718
rect 303804 326392 303856 326398
rect 303804 326334 303856 326340
rect 303620 326324 303672 326330
rect 303620 326266 303672 326272
rect 303908 321502 303936 340068
rect 304000 340054 304198 340082
rect 304276 340054 304474 340082
rect 304552 340054 304658 340082
rect 304736 340054 304934 340082
rect 304000 335782 304028 340054
rect 303988 335776 304040 335782
rect 303988 335718 304040 335724
rect 303988 335640 304040 335646
rect 304276 335594 304304 340054
rect 304552 335646 304580 340054
rect 303988 335582 304040 335588
rect 304000 326346 304028 335582
rect 304092 335566 304304 335594
rect 304540 335640 304592 335646
rect 304540 335582 304592 335588
rect 304092 326466 304120 335566
rect 304736 331294 304764 340054
rect 304724 331288 304776 331294
rect 304724 331230 304776 331236
rect 304264 331220 304316 331226
rect 304264 331162 304316 331168
rect 304276 326482 304304 331162
rect 305000 329996 305052 330002
rect 305000 329938 305052 329944
rect 304080 326460 304132 326466
rect 304276 326454 304764 326482
rect 304080 326402 304132 326408
rect 304632 326392 304684 326398
rect 304000 326318 304580 326346
rect 304632 326334 304684 326340
rect 303896 321496 303948 321502
rect 303896 321438 303948 321444
rect 304448 321496 304500 321502
rect 304448 321438 304500 321444
rect 304460 17406 304488 321438
rect 304448 17400 304500 17406
rect 304448 17342 304500 17348
rect 304552 17338 304580 326318
rect 304644 17474 304672 326334
rect 304632 17468 304684 17474
rect 304632 17410 304684 17416
rect 304540 17332 304592 17338
rect 304540 17274 304592 17280
rect 304736 17270 304764 326454
rect 304816 326460 304868 326466
rect 304816 326402 304868 326408
rect 304828 18086 304856 326402
rect 305012 326330 305040 329938
rect 305104 326398 305132 340068
rect 305196 336977 305224 340190
rect 317972 340138 318024 340144
rect 318444 340190 318642 340218
rect 305656 338042 305684 340068
rect 305472 338014 305684 338042
rect 305748 340054 305854 340082
rect 306024 340054 306130 340082
rect 306406 340054 306512 340082
rect 305182 336968 305238 336977
rect 305182 336903 305238 336912
rect 305366 336832 305422 336841
rect 305366 336767 305422 336776
rect 305380 336734 305408 336767
rect 305368 336728 305420 336734
rect 305368 336670 305420 336676
rect 305184 335640 305236 335646
rect 305184 335582 305236 335588
rect 305196 326466 305224 335582
rect 305472 330002 305500 338014
rect 305552 336728 305604 336734
rect 305552 336670 305604 336676
rect 305460 329996 305512 330002
rect 305460 329938 305512 329944
rect 305564 328386 305592 336670
rect 305748 335646 305776 340054
rect 305736 335640 305788 335646
rect 305736 335582 305788 335588
rect 305472 328358 305592 328386
rect 305184 326460 305236 326466
rect 305184 326402 305236 326408
rect 305092 326392 305144 326398
rect 305092 326334 305144 326340
rect 304908 326324 304960 326330
rect 304908 326266 304960 326272
rect 305000 326324 305052 326330
rect 305000 326266 305052 326272
rect 304816 18080 304868 18086
rect 304816 18022 304868 18028
rect 304920 18018 304948 326266
rect 305472 323610 305500 328358
rect 305460 323604 305512 323610
rect 305460 323546 305512 323552
rect 305920 323604 305972 323610
rect 305920 323546 305972 323552
rect 304908 18012 304960 18018
rect 304908 17954 304960 17960
rect 305932 17785 305960 323546
rect 305918 17776 305974 17785
rect 305918 17711 305974 17720
rect 304724 17264 304776 17270
rect 304724 17206 304776 17212
rect 304644 15286 304856 15314
rect 304644 15230 304672 15286
rect 304632 15224 304684 15230
rect 304632 15166 304684 15172
rect 303528 8152 303580 8158
rect 303528 8094 303580 8100
rect 304828 8022 304856 15286
rect 304908 15224 304960 15230
rect 304908 15166 304960 15172
rect 304920 8090 304948 15166
rect 306024 11286 306052 340054
rect 306484 326466 306512 340054
rect 306196 326460 306248 326466
rect 306196 326402 306248 326408
rect 306472 326460 306524 326466
rect 306472 326402 306524 326408
rect 306104 326392 306156 326398
rect 306104 326334 306156 326340
rect 306012 11280 306064 11286
rect 306012 11222 306064 11228
rect 304908 8084 304960 8090
rect 304908 8026 304960 8032
rect 304816 8016 304868 8022
rect 304816 7958 304868 7964
rect 306116 7954 306144 326334
rect 306104 7948 306156 7954
rect 306104 7890 306156 7896
rect 306208 7886 306236 326402
rect 306576 326398 306604 340068
rect 306656 335640 306708 335646
rect 306656 335582 306708 335588
rect 306668 328574 306696 335582
rect 306748 333328 306800 333334
rect 306748 333270 306800 333276
rect 306656 328568 306708 328574
rect 306656 328510 306708 328516
rect 306564 326392 306616 326398
rect 306564 326334 306616 326340
rect 306288 326324 306340 326330
rect 306288 326266 306340 326272
rect 306196 7880 306248 7886
rect 306196 7822 306248 7828
rect 303804 7744 303856 7750
rect 303804 7686 303856 7692
rect 300768 7540 300820 7546
rect 300768 7482 300820 7488
rect 300676 7472 300728 7478
rect 300676 7414 300728 7420
rect 301412 5160 301464 5166
rect 301412 5102 301464 5108
rect 301424 480 301452 5102
rect 302608 5092 302660 5098
rect 302608 5034 302660 5040
rect 302620 480 302648 5034
rect 303816 480 303844 7686
rect 305000 5024 305052 5030
rect 305000 4966 305052 4972
rect 305012 480 305040 4966
rect 306196 4956 306248 4962
rect 306196 4898 306248 4904
rect 306208 480 306236 4898
rect 306300 4282 306328 326266
rect 306760 316418 306788 333270
rect 306852 316690 306880 340068
rect 306944 340054 307142 340082
rect 307326 340054 307432 340082
rect 306944 335646 306972 340054
rect 306932 335640 306984 335646
rect 306932 335582 306984 335588
rect 306852 316662 307340 316690
rect 306760 316390 307248 316418
rect 307220 15230 307248 316390
rect 307208 15224 307260 15230
rect 307208 15166 307260 15172
rect 307312 12442 307340 316662
rect 307024 12436 307076 12442
rect 307024 12378 307076 12384
rect 307300 12436 307352 12442
rect 307300 12378 307352 12384
rect 307036 11354 307064 12378
rect 307024 11348 307076 11354
rect 307024 11290 307076 11296
rect 307404 7818 307432 340054
rect 307496 340054 307602 340082
rect 307496 333334 307524 340054
rect 307760 335708 307812 335714
rect 307760 335650 307812 335656
rect 307484 333328 307536 333334
rect 307484 333270 307536 333276
rect 307576 328568 307628 328574
rect 307576 328510 307628 328516
rect 307484 326392 307536 326398
rect 307484 326334 307536 326340
rect 307496 7818 307524 326334
rect 307392 7812 307444 7818
rect 307392 7754 307444 7760
rect 307484 7812 307536 7818
rect 307484 7754 307536 7760
rect 307392 7676 307444 7682
rect 307392 7618 307444 7624
rect 306288 4276 306340 4282
rect 306288 4218 306340 4224
rect 307404 480 307432 7618
rect 307588 4418 307616 328510
rect 307668 326460 307720 326466
rect 307668 326402 307720 326408
rect 307576 4412 307628 4418
rect 307576 4354 307628 4360
rect 307680 4350 307708 326402
rect 307772 326262 307800 335650
rect 307864 326534 307892 340068
rect 307944 335640 307996 335646
rect 307944 335582 307996 335588
rect 307852 326528 307904 326534
rect 307852 326470 307904 326476
rect 307956 326330 307984 335582
rect 308048 326466 308076 340068
rect 308338 340054 308536 340082
rect 308508 335594 308536 340054
rect 308600 335714 308628 340068
rect 308692 340054 308798 340082
rect 308876 340054 309074 340082
rect 309244 340054 309350 340082
rect 308588 335708 308640 335714
rect 308588 335650 308640 335656
rect 308692 335646 308720 340054
rect 308680 335640 308732 335646
rect 308508 335566 308628 335594
rect 308680 335582 308732 335588
rect 308128 332988 308180 332994
rect 308128 332930 308180 332936
rect 308036 326460 308088 326466
rect 308036 326402 308088 326408
rect 308140 326398 308168 332930
rect 308128 326392 308180 326398
rect 308128 326334 308180 326340
rect 307944 326324 307996 326330
rect 307944 326266 307996 326272
rect 307760 326256 307812 326262
rect 307760 326198 307812 326204
rect 308402 16280 308458 16289
rect 308402 16215 308458 16224
rect 308416 15609 308444 16215
rect 308402 15600 308458 15609
rect 308402 15535 308458 15544
rect 308600 12442 308628 335566
rect 308876 332994 308904 340054
rect 309140 338972 309192 338978
rect 309140 338914 309192 338920
rect 308864 332988 308916 332994
rect 308864 332930 308916 332936
rect 308956 326528 309008 326534
rect 308956 326470 309008 326476
rect 308864 326460 308916 326466
rect 308864 326402 308916 326408
rect 308680 326392 308732 326398
rect 308680 326334 308732 326340
rect 308496 12436 308548 12442
rect 308496 12378 308548 12384
rect 308588 12436 308640 12442
rect 308588 12378 308640 12384
rect 308508 11490 308536 12378
rect 308692 11558 308720 326334
rect 308772 326324 308824 326330
rect 308772 326266 308824 326272
rect 308680 11552 308732 11558
rect 308680 11494 308732 11500
rect 308496 11484 308548 11490
rect 308496 11426 308548 11432
rect 308784 8265 308812 326266
rect 308770 8256 308826 8265
rect 308770 8191 308826 8200
rect 308876 7682 308904 326402
rect 308864 7676 308916 7682
rect 308864 7618 308916 7624
rect 308588 4888 308640 4894
rect 308588 4830 308640 4836
rect 307668 4344 307720 4350
rect 307668 4286 307720 4292
rect 308600 480 308628 4830
rect 308968 4486 308996 326470
rect 309152 326466 309180 338914
rect 309140 326460 309192 326466
rect 309140 326402 309192 326408
rect 309244 326330 309272 340054
rect 309520 338978 309548 340068
rect 309612 340054 309810 340082
rect 309508 338972 309560 338978
rect 309508 338914 309560 338920
rect 309612 335594 309640 340054
rect 310072 338162 310100 340068
rect 310164 340054 310270 340082
rect 309876 338156 309928 338162
rect 309876 338098 309928 338104
rect 310060 338156 310112 338162
rect 310060 338098 310112 338104
rect 309428 335566 309640 335594
rect 309232 326324 309284 326330
rect 309232 326266 309284 326272
rect 309048 326256 309100 326262
rect 309048 326198 309100 326204
rect 309060 4554 309088 326198
rect 309428 321570 309456 335566
rect 309888 331294 309916 338098
rect 309876 331288 309928 331294
rect 309876 331230 309928 331236
rect 309692 331220 309744 331226
rect 309692 331162 309744 331168
rect 309704 328386 309732 331162
rect 309520 328358 309732 328386
rect 309520 323610 309548 328358
rect 309508 323604 309560 323610
rect 309508 323546 309560 323552
rect 309416 321564 309468 321570
rect 309416 321506 309468 321512
rect 310060 321564 310112 321570
rect 310060 321506 310112 321512
rect 310072 309942 310100 321506
rect 310060 309936 310112 309942
rect 310060 309878 310112 309884
rect 310060 309800 310112 309806
rect 310060 309742 310112 309748
rect 310072 12442 310100 309742
rect 309968 12436 310020 12442
rect 309968 12378 310020 12384
rect 310060 12436 310112 12442
rect 310060 12378 310112 12384
rect 309980 11626 310008 12378
rect 309968 11620 310020 11626
rect 309968 11562 310020 11568
rect 310164 7993 310192 340054
rect 310532 335646 310560 340068
rect 310624 340054 310822 340082
rect 310520 335640 310572 335646
rect 310520 335582 310572 335588
rect 310244 326460 310296 326466
rect 310244 326402 310296 326408
rect 310256 8129 310284 326402
rect 310624 326398 310652 340054
rect 310992 335714 311020 340068
rect 311084 340054 311282 340082
rect 310980 335708 311032 335714
rect 310980 335650 311032 335656
rect 310704 335640 310756 335646
rect 311084 335594 311112 340054
rect 311544 338042 311572 340068
rect 310704 335582 310756 335588
rect 310612 326392 310664 326398
rect 310612 326334 310664 326340
rect 310428 326324 310480 326330
rect 310428 326266 310480 326272
rect 310336 323604 310388 323610
rect 310336 323546 310388 323552
rect 310242 8120 310298 8129
rect 310242 8055 310298 8064
rect 310150 7984 310206 7993
rect 310150 7919 310206 7928
rect 309782 5536 309838 5545
rect 309782 5471 309838 5480
rect 309048 4548 309100 4554
rect 309048 4490 309100 4496
rect 308956 4480 309008 4486
rect 308956 4422 309008 4428
rect 309796 480 309824 5471
rect 310348 4690 310376 323546
rect 310336 4684 310388 4690
rect 310336 4626 310388 4632
rect 310440 4622 310468 326266
rect 310716 326262 310744 335582
rect 310900 335566 311112 335594
rect 311452 338014 311572 338042
rect 311636 340054 311742 340082
rect 310704 326256 310756 326262
rect 310704 326198 310756 326204
rect 310900 321570 310928 335566
rect 311072 335504 311124 335510
rect 311072 335446 311124 335452
rect 311084 326346 311112 335446
rect 311452 331906 311480 338014
rect 311636 335510 311664 340054
rect 312004 335850 312032 340068
rect 312096 340054 312294 340082
rect 312372 340054 312478 340082
rect 312648 340054 312754 340082
rect 313030 340054 313136 340082
rect 311992 335844 312044 335850
rect 311992 335786 312044 335792
rect 311716 335708 311768 335714
rect 312096 335696 312124 340054
rect 311716 335650 311768 335656
rect 311912 335668 312124 335696
rect 311624 335504 311676 335510
rect 311624 335446 311676 335452
rect 311256 331900 311308 331906
rect 311256 331842 311308 331848
rect 311440 331900 311492 331906
rect 311440 331842 311492 331848
rect 311268 326466 311296 331842
rect 311728 326618 311756 335650
rect 311636 326590 311756 326618
rect 311256 326460 311308 326466
rect 311256 326402 311308 326408
rect 311084 326318 311572 326346
rect 311440 326256 311492 326262
rect 311440 326198 311492 326204
rect 310888 321564 310940 321570
rect 310888 321506 310940 321512
rect 311348 321564 311400 321570
rect 311348 321506 311400 321512
rect 311360 309942 311388 321506
rect 311348 309936 311400 309942
rect 311348 309878 311400 309884
rect 311348 309800 311400 309806
rect 311348 309742 311400 309748
rect 311360 12374 311388 309742
rect 311348 12368 311400 12374
rect 311348 12310 311400 12316
rect 311452 11694 311480 326198
rect 311440 11688 311492 11694
rect 311440 11630 311492 11636
rect 311544 7857 311572 326318
rect 311530 7848 311586 7857
rect 311530 7783 311586 7792
rect 311636 7614 311664 326590
rect 311912 326534 311940 335668
rect 312176 335640 312228 335646
rect 312176 335582 312228 335588
rect 312084 335572 312136 335578
rect 312084 335514 312136 335520
rect 311900 326528 311952 326534
rect 311900 326470 311952 326476
rect 312096 326466 312124 335514
rect 311716 326460 311768 326466
rect 311716 326402 311768 326408
rect 312084 326460 312136 326466
rect 312084 326402 312136 326408
rect 310980 7608 311032 7614
rect 310980 7550 311032 7556
rect 311624 7608 311676 7614
rect 311624 7550 311676 7556
rect 310428 4616 310480 4622
rect 310428 4558 310480 4564
rect 310992 480 311020 7550
rect 311728 5506 311756 326402
rect 311808 326392 311860 326398
rect 311808 326334 311860 326340
rect 311716 5500 311768 5506
rect 311716 5442 311768 5448
rect 311820 4758 311848 326334
rect 312188 326330 312216 335582
rect 312372 326398 312400 340054
rect 312544 335844 312596 335850
rect 312544 335786 312596 335792
rect 312360 326392 312412 326398
rect 312360 326334 312412 326340
rect 312176 326324 312228 326330
rect 312176 326266 312228 326272
rect 312556 311794 312584 335786
rect 312648 335578 312676 340054
rect 312636 335572 312688 335578
rect 312636 335514 312688 335520
rect 313108 335492 313136 340054
rect 313200 335646 313228 340068
rect 313490 340054 313596 340082
rect 313372 336048 313424 336054
rect 313372 335990 313424 335996
rect 313188 335640 313240 335646
rect 313188 335582 313240 335588
rect 313280 335640 313332 335646
rect 313280 335582 313332 335588
rect 313108 335464 313228 335492
rect 313096 326528 313148 326534
rect 313096 326470 313148 326476
rect 312820 326460 312872 326466
rect 312820 326402 312872 326408
rect 312556 311766 312768 311794
rect 311990 16824 312046 16833
rect 311990 16759 312046 16768
rect 311898 16688 311954 16697
rect 312004 16674 312032 16759
rect 311954 16646 312032 16674
rect 311898 16623 311954 16632
rect 312740 12374 312768 311766
rect 312728 12368 312780 12374
rect 312728 12310 312780 12316
rect 312832 12306 312860 326402
rect 312912 326392 312964 326398
rect 312912 326334 312964 326340
rect 312820 12300 312872 12306
rect 312820 12242 312872 12248
rect 312924 7721 312952 326334
rect 313004 326324 313056 326330
rect 313004 326266 313056 326272
rect 312910 7712 312966 7721
rect 312910 7647 312966 7656
rect 313016 7585 313044 326266
rect 313002 7576 313058 7585
rect 313002 7511 313058 7520
rect 313108 5438 313136 326470
rect 313096 5432 313148 5438
rect 313096 5374 313148 5380
rect 313200 5370 313228 335464
rect 313292 326534 313320 335582
rect 313280 326528 313332 326534
rect 313280 326470 313332 326476
rect 313384 326330 313412 335990
rect 313568 335986 313596 340054
rect 313660 340054 313766 340082
rect 313950 340054 314148 340082
rect 313660 336054 313688 340054
rect 313648 336048 313700 336054
rect 313648 335990 313700 335996
rect 313556 335980 313608 335986
rect 313556 335922 313608 335928
rect 313556 335776 313608 335782
rect 313556 335718 313608 335724
rect 313568 326466 313596 335718
rect 313648 335708 313700 335714
rect 313648 335650 313700 335656
rect 313556 326460 313608 326466
rect 313556 326402 313608 326408
rect 313660 326398 313688 335650
rect 314120 331922 314148 340054
rect 314212 335714 314240 340068
rect 314304 340054 314502 340082
rect 314686 340054 314884 340082
rect 314962 340054 315160 340082
rect 314200 335708 314252 335714
rect 314200 335650 314252 335656
rect 314304 335646 314332 340054
rect 314752 335708 314804 335714
rect 314752 335650 314804 335656
rect 314292 335640 314344 335646
rect 314292 335582 314344 335588
rect 314120 331894 314240 331922
rect 313648 326392 313700 326398
rect 313648 326334 313700 326340
rect 313372 326324 313424 326330
rect 313372 326266 313424 326272
rect 314212 143478 314240 331894
rect 314568 326528 314620 326534
rect 314568 326470 314620 326476
rect 314384 326460 314436 326466
rect 314384 326402 314436 326408
rect 314292 326392 314344 326398
rect 314292 326334 314344 326340
rect 314304 143546 314332 326334
rect 314396 143546 314424 326402
rect 314476 326324 314528 326330
rect 314476 326266 314528 326272
rect 314292 143540 314344 143546
rect 314292 143482 314344 143488
rect 314384 143540 314436 143546
rect 314384 143482 314436 143488
rect 314200 143472 314252 143478
rect 314200 143414 314252 143420
rect 314292 143404 314344 143410
rect 314292 143346 314344 143352
rect 314200 143336 314252 143342
rect 314200 143278 314252 143284
rect 314212 77246 314240 143278
rect 314200 77240 314252 77246
rect 314200 77182 314252 77188
rect 314200 67652 314252 67658
rect 314200 67594 314252 67600
rect 314212 66230 314240 67594
rect 314200 66224 314252 66230
rect 314200 66166 314252 66172
rect 314200 56636 314252 56642
rect 314200 56578 314252 56584
rect 314212 46918 314240 56578
rect 314200 46912 314252 46918
rect 314200 46854 314252 46860
rect 314200 37324 314252 37330
rect 314200 37266 314252 37272
rect 314212 27606 314240 37266
rect 314200 27600 314252 27606
rect 314200 27542 314252 27548
rect 314200 18012 314252 18018
rect 314200 17954 314252 17960
rect 314212 17649 314240 17954
rect 314198 17640 314254 17649
rect 314198 17575 314254 17584
rect 314304 12170 314332 143346
rect 314384 138508 314436 138514
rect 314384 138450 314436 138456
rect 314396 124098 314424 138450
rect 314384 124092 314436 124098
rect 314384 124034 314436 124040
rect 314384 123956 314436 123962
rect 314384 123898 314436 123904
rect 314396 77178 314424 123898
rect 314384 77172 314436 77178
rect 314384 77114 314436 77120
rect 314384 77036 314436 77042
rect 314384 76978 314436 76984
rect 314396 12238 314424 76978
rect 314384 12232 314436 12238
rect 314384 12174 314436 12180
rect 314292 12164 314344 12170
rect 314292 12106 314344 12112
rect 314384 11076 314436 11082
rect 314384 11018 314436 11024
rect 313370 5400 313426 5409
rect 313188 5364 313240 5370
rect 313370 5335 313426 5344
rect 313188 5306 313240 5312
rect 312176 4820 312228 4826
rect 312176 4762 312228 4768
rect 311808 4752 311860 4758
rect 311808 4694 311860 4700
rect 311806 4176 311862 4185
rect 311806 4111 311862 4120
rect 311820 3670 311848 4111
rect 311808 3664 311860 3670
rect 311808 3606 311860 3612
rect 312188 480 312216 4762
rect 313384 480 313412 5335
rect 314396 5234 314424 11018
rect 314488 5302 314516 326266
rect 314580 11082 314608 326470
rect 314764 326398 314792 335650
rect 314752 326392 314804 326398
rect 314752 326334 314804 326340
rect 314856 326262 314884 340054
rect 315028 335504 315080 335510
rect 315028 335446 315080 335452
rect 314844 326256 314896 326262
rect 314844 326198 314896 326204
rect 315040 318782 315068 335446
rect 315132 326380 315160 340054
rect 315224 326534 315252 340068
rect 315316 340054 315422 340082
rect 315698 340054 315804 340082
rect 315316 335510 315344 340054
rect 315304 335504 315356 335510
rect 315304 335446 315356 335452
rect 315212 326528 315264 326534
rect 315212 326470 315264 326476
rect 315132 326352 315712 326380
rect 315580 326256 315632 326262
rect 315580 326198 315632 326204
rect 315028 318776 315080 318782
rect 315028 318718 315080 318724
rect 315488 318776 315540 318782
rect 315488 318718 315540 318724
rect 315500 17377 315528 318718
rect 315592 17513 315620 326198
rect 315578 17504 315634 17513
rect 315578 17439 315634 17448
rect 315486 17368 315542 17377
rect 315486 17303 315542 17312
rect 315684 12102 315712 326352
rect 315672 12096 315724 12102
rect 315672 12038 315724 12044
rect 315776 12034 315804 340054
rect 315868 340054 315974 340082
rect 316158 340054 316264 340082
rect 315868 335714 315896 340054
rect 315856 335708 315908 335714
rect 315856 335650 315908 335656
rect 316132 335640 316184 335646
rect 316132 335582 316184 335588
rect 315856 326528 315908 326534
rect 315856 326470 315908 326476
rect 315764 12028 315816 12034
rect 315764 11970 315816 11976
rect 314568 11076 314620 11082
rect 314568 11018 314620 11024
rect 314568 9172 314620 9178
rect 314568 9114 314620 9120
rect 314476 5296 314528 5302
rect 314476 5238 314528 5244
rect 314384 5228 314436 5234
rect 314384 5170 314436 5176
rect 313922 4176 313978 4185
rect 313922 4111 313978 4120
rect 313936 3670 313964 4111
rect 313924 3664 313976 3670
rect 313924 3606 313976 3612
rect 314580 480 314608 9114
rect 315868 5166 315896 326470
rect 315948 326392 316000 326398
rect 315948 326334 316000 326340
rect 315856 5160 315908 5166
rect 315762 5128 315818 5137
rect 315856 5102 315908 5108
rect 315960 5098 315988 326334
rect 316144 316606 316172 335582
rect 316236 326398 316264 340054
rect 316328 340054 316434 340082
rect 316604 340054 316710 340082
rect 316224 326392 316276 326398
rect 316224 326334 316276 326340
rect 316328 326244 316356 340054
rect 316500 338972 316552 338978
rect 316500 338914 316552 338920
rect 316512 326380 316540 338914
rect 316604 326482 316632 340054
rect 316880 338978 316908 340068
rect 316972 340054 317170 340082
rect 317446 340054 317552 340082
rect 317630 340054 317828 340082
rect 316868 338972 316920 338978
rect 316868 338914 316920 338920
rect 316972 335646 317000 340054
rect 316960 335640 317012 335646
rect 316960 335582 317012 335588
rect 317524 330342 317552 340054
rect 317696 335844 317748 335850
rect 317696 335786 317748 335792
rect 317512 330336 317564 330342
rect 317512 330278 317564 330284
rect 316604 326454 317368 326482
rect 317236 326392 317288 326398
rect 316512 326352 317184 326380
rect 316328 326216 317092 326244
rect 316132 316600 316184 316606
rect 316132 316542 316184 316548
rect 316868 316600 316920 316606
rect 316868 316542 316920 316548
rect 316880 307766 316908 316542
rect 316868 307760 316920 307766
rect 316868 307702 316920 307708
rect 316960 298172 317012 298178
rect 316960 298114 317012 298120
rect 316972 114510 317000 298114
rect 316960 114504 317012 114510
rect 316960 114446 317012 114452
rect 316960 104916 317012 104922
rect 316960 104858 317012 104864
rect 316972 67658 317000 104858
rect 317064 77246 317092 326216
rect 317156 124166 317184 326352
rect 317236 326334 317288 326340
rect 317144 124160 317196 124166
rect 317144 124102 317196 124108
rect 317144 117564 317196 117570
rect 317144 117506 317196 117512
rect 317156 114510 317184 117506
rect 317144 114504 317196 114510
rect 317144 114446 317196 114452
rect 317248 114442 317276 326334
rect 317340 124166 317368 326454
rect 317708 326330 317736 335786
rect 317800 335578 317828 340054
rect 317984 340054 318182 340082
rect 318260 340054 318366 340082
rect 317880 338156 317932 338162
rect 317880 338098 317932 338104
rect 317788 335572 317840 335578
rect 317788 335514 317840 335520
rect 317696 326324 317748 326330
rect 317696 326266 317748 326272
rect 317892 315246 317920 338098
rect 317984 335850 318012 340054
rect 317972 335844 318024 335850
rect 317972 335786 318024 335792
rect 318260 335696 318288 340054
rect 317984 335668 318288 335696
rect 317984 326466 318012 335668
rect 318064 335572 318116 335578
rect 318064 335514 318116 335520
rect 317972 326460 318024 326466
rect 317972 326402 318024 326408
rect 318076 326398 318104 335514
rect 318444 335345 318472 340190
rect 318812 340054 318918 340082
rect 318154 335336 318210 335345
rect 318154 335271 318210 335280
rect 318430 335336 318486 335345
rect 318430 335271 318486 335280
rect 318064 326392 318116 326398
rect 318064 326334 318116 326340
rect 318168 325718 318196 335271
rect 318616 330336 318668 330342
rect 318616 330278 318668 330284
rect 318432 326460 318484 326466
rect 318432 326402 318484 326408
rect 318156 325712 318208 325718
rect 318156 325654 318208 325660
rect 318248 325712 318300 325718
rect 318248 325654 318300 325660
rect 318260 322266 318288 325654
rect 318076 322238 318288 322266
rect 317880 315240 317932 315246
rect 317880 315182 317932 315188
rect 318076 307086 318104 322238
rect 318248 315240 318300 315246
rect 318248 315182 318300 315188
rect 318064 307080 318116 307086
rect 318064 307022 318116 307028
rect 317328 124160 317380 124166
rect 317328 124102 317380 124108
rect 317328 115592 317380 115598
rect 317328 115534 317380 115540
rect 317340 114510 317368 115534
rect 317328 114504 317380 114510
rect 317328 114446 317380 114452
rect 317236 114436 317288 114442
rect 317236 114378 317288 114384
rect 317328 109744 317380 109750
rect 317328 109686 317380 109692
rect 317144 107636 317196 107642
rect 317144 107578 317196 107584
rect 317052 77240 317104 77246
rect 317052 77182 317104 77188
rect 317052 77104 317104 77110
rect 317052 77046 317104 77052
rect 316868 67652 316920 67658
rect 316868 67594 316920 67600
rect 316960 67652 317012 67658
rect 316960 67594 317012 67600
rect 316880 11898 316908 67594
rect 317064 11966 317092 77046
rect 317052 11960 317104 11966
rect 317052 11902 317104 11908
rect 316868 11892 316920 11898
rect 316868 11834 316920 11840
rect 317156 9489 317184 107578
rect 317236 106140 317288 106146
rect 317236 106082 317288 106088
rect 317142 9480 317198 9489
rect 317142 9415 317198 9424
rect 317248 9110 317276 106082
rect 317236 9104 317288 9110
rect 317236 9046 317288 9052
rect 317050 5264 317106 5273
rect 317050 5199 317106 5208
rect 315762 5063 315818 5072
rect 315948 5092 316000 5098
rect 315776 480 315804 5063
rect 315948 5034 316000 5040
rect 316604 3738 317000 3754
rect 316604 3732 317012 3738
rect 316604 3726 316960 3732
rect 316604 3670 316632 3726
rect 316960 3674 317012 3680
rect 316592 3664 316644 3670
rect 317064 3618 317092 5199
rect 317340 5030 317368 109686
rect 318260 77246 318288 315182
rect 318340 307080 318392 307086
rect 318340 307022 318392 307028
rect 318248 77240 318300 77246
rect 318248 77182 318300 77188
rect 318156 67652 318208 67658
rect 318156 67594 318208 67600
rect 318168 11830 318196 67594
rect 318156 11824 318208 11830
rect 318156 11766 318208 11772
rect 318352 11762 318380 307022
rect 318340 11756 318392 11762
rect 318340 11698 318392 11704
rect 318444 9353 318472 326402
rect 318524 326392 318576 326398
rect 318524 326334 318576 326340
rect 318430 9344 318486 9353
rect 318430 9279 318486 9288
rect 318536 9178 318564 326334
rect 318064 9172 318116 9178
rect 318064 9114 318116 9120
rect 318524 9172 318576 9178
rect 318524 9114 318576 9120
rect 317328 5024 317380 5030
rect 317328 4966 317380 4972
rect 316592 3606 316644 3612
rect 316972 3590 317092 3618
rect 316972 480 317000 3590
rect 318076 480 318104 9114
rect 318628 4962 318656 330278
rect 318812 326534 318840 340054
rect 318984 335640 319036 335646
rect 318984 335582 319036 335588
rect 318800 326528 318852 326534
rect 318800 326470 318852 326476
rect 318996 326330 319024 335582
rect 319088 326466 319116 340068
rect 319180 340054 319378 340082
rect 319456 340054 319654 340082
rect 319838 340054 319944 340082
rect 319076 326460 319128 326466
rect 319076 326402 319128 326408
rect 319180 326398 319208 340054
rect 319456 335646 319484 340054
rect 319536 338156 319588 338162
rect 319536 338098 319588 338104
rect 319444 335640 319496 335646
rect 319444 335582 319496 335588
rect 319548 335322 319576 338098
rect 319456 335294 319576 335322
rect 319456 328438 319484 335294
rect 319444 328432 319496 328438
rect 319444 328374 319496 328380
rect 319812 326460 319864 326466
rect 319812 326402 319864 326408
rect 319168 326392 319220 326398
rect 319168 326334 319220 326340
rect 319720 326392 319772 326398
rect 319720 326334 319772 326340
rect 318708 326324 318760 326330
rect 318708 326266 318760 326272
rect 318984 326324 319036 326330
rect 318984 326266 319036 326272
rect 318616 4956 318668 4962
rect 318616 4898 318668 4904
rect 318720 4894 318748 326266
rect 319444 325712 319496 325718
rect 319442 325680 319444 325689
rect 319496 325680 319498 325689
rect 319442 325615 319498 325624
rect 319626 325680 319682 325689
rect 319626 325615 319682 325624
rect 319640 316130 319668 325615
rect 319444 316124 319496 316130
rect 319444 316066 319496 316072
rect 319628 316124 319680 316130
rect 319628 316066 319680 316072
rect 319456 315994 319484 316066
rect 319444 315988 319496 315994
rect 319444 315930 319496 315936
rect 319628 306400 319680 306406
rect 319628 306342 319680 306348
rect 319640 298110 319668 306342
rect 319628 298104 319680 298110
rect 319628 298046 319680 298052
rect 319628 287088 319680 287094
rect 319628 287030 319680 287036
rect 319640 277409 319668 287030
rect 319442 277400 319498 277409
rect 319442 277335 319498 277344
rect 319626 277400 319682 277409
rect 319626 277335 319682 277344
rect 319456 267782 319484 277335
rect 319444 267776 319496 267782
rect 319444 267718 319496 267724
rect 319628 267776 319680 267782
rect 319628 267718 319680 267724
rect 319640 258058 319668 267718
rect 319628 258052 319680 258058
rect 319628 257994 319680 258000
rect 319628 240168 319680 240174
rect 319628 240110 319680 240116
rect 319640 238746 319668 240110
rect 319444 238740 319496 238746
rect 319444 238682 319496 238688
rect 319628 238740 319680 238746
rect 319628 238682 319680 238688
rect 319456 229129 319484 238682
rect 319442 229120 319498 229129
rect 319442 229055 319498 229064
rect 319626 229120 319682 229129
rect 319626 229055 319682 229064
rect 319640 219434 319668 229055
rect 319628 219428 319680 219434
rect 319628 219370 319680 219376
rect 319628 209840 319680 209846
rect 319628 209782 319680 209788
rect 319640 200122 319668 209782
rect 319628 200116 319680 200122
rect 319628 200058 319680 200064
rect 319628 190528 319680 190534
rect 319628 190470 319680 190476
rect 319640 180810 319668 190470
rect 319628 180804 319680 180810
rect 319628 180746 319680 180752
rect 319628 171148 319680 171154
rect 319628 171090 319680 171096
rect 319640 161430 319668 171090
rect 319628 161424 319680 161430
rect 319628 161366 319680 161372
rect 319628 151836 319680 151842
rect 319628 151778 319680 151784
rect 319640 143721 319668 151778
rect 319626 143712 319682 143721
rect 319626 143647 319682 143656
rect 319626 143576 319682 143585
rect 319626 143511 319682 143520
rect 319640 142118 319668 143511
rect 319628 142112 319680 142118
rect 319628 142054 319680 142060
rect 319628 132524 319680 132530
rect 319628 132466 319680 132472
rect 319640 122806 319668 132466
rect 319628 122800 319680 122806
rect 319628 122742 319680 122748
rect 319628 113212 319680 113218
rect 319628 113154 319680 113160
rect 319640 103494 319668 113154
rect 319628 103488 319680 103494
rect 319628 103430 319680 103436
rect 319628 93900 319680 93906
rect 319628 93842 319680 93848
rect 319640 84182 319668 93842
rect 319628 84176 319680 84182
rect 319628 84118 319680 84124
rect 319628 74588 319680 74594
rect 319628 74530 319680 74536
rect 319640 64870 319668 74530
rect 319628 64864 319680 64870
rect 319628 64806 319680 64812
rect 319628 46980 319680 46986
rect 319628 46922 319680 46928
rect 319640 45558 319668 46922
rect 319628 45552 319680 45558
rect 319628 45494 319680 45500
rect 319628 35964 319680 35970
rect 319628 35906 319680 35912
rect 319640 31822 319668 35906
rect 319628 31816 319680 31822
rect 319628 31758 319680 31764
rect 319536 31748 319588 31754
rect 319536 31690 319588 31696
rect 319548 12209 319576 31690
rect 319732 12345 319760 326334
rect 319718 12336 319774 12345
rect 319718 12271 319774 12280
rect 319534 12200 319590 12209
rect 319534 12135 319590 12144
rect 319824 9217 319852 326402
rect 319810 9208 319866 9217
rect 319810 9143 319866 9152
rect 319916 9081 319944 340054
rect 320100 338162 320128 340068
rect 320298 340054 320404 340082
rect 320088 338156 320140 338162
rect 320088 338098 320140 338104
rect 320180 335980 320232 335986
rect 320180 335922 320232 335928
rect 320192 335238 320220 335922
rect 320180 335232 320232 335238
rect 320180 335174 320232 335180
rect 320376 330614 320404 340054
rect 320468 340054 320574 340082
rect 320364 330608 320416 330614
rect 320364 330550 320416 330556
rect 320088 326528 320140 326534
rect 320088 326470 320140 326476
rect 319996 326324 320048 326330
rect 319996 326266 320048 326272
rect 319902 9072 319958 9081
rect 319902 9007 319958 9016
rect 320008 5545 320036 326266
rect 319994 5536 320050 5545
rect 319994 5471 320050 5480
rect 319258 4992 319314 5001
rect 319258 4927 319314 4936
rect 318708 4888 318760 4894
rect 318708 4830 318760 4836
rect 319272 480 319300 4927
rect 320100 4826 320128 326470
rect 320468 326398 320496 340054
rect 320836 335986 320864 340068
rect 320928 340054 321034 340082
rect 321112 340054 321310 340082
rect 320824 335980 320876 335986
rect 320824 335922 320876 335928
rect 320640 335640 320692 335646
rect 320640 335582 320692 335588
rect 320456 326392 320508 326398
rect 320652 326380 320680 335582
rect 320928 335442 320956 340054
rect 321112 335646 321140 340054
rect 321100 335640 321152 335646
rect 321100 335582 321152 335588
rect 320916 335436 320968 335442
rect 320916 335378 320968 335384
rect 321468 335436 321520 335442
rect 321468 335378 321520 335384
rect 321376 330608 321428 330614
rect 321376 330550 321428 330556
rect 321284 326392 321336 326398
rect 320652 326352 321232 326380
rect 320456 326334 320508 326340
rect 320272 325712 320324 325718
rect 320272 325654 320324 325660
rect 320284 315994 320312 325654
rect 320272 315988 320324 315994
rect 320272 315930 320324 315936
rect 321100 306400 321152 306406
rect 321100 306342 321152 306348
rect 321112 298110 321140 306342
rect 321100 298104 321152 298110
rect 321100 298046 321152 298052
rect 321100 288516 321152 288522
rect 321100 288458 321152 288464
rect 321112 278769 321140 288458
rect 320914 278760 320970 278769
rect 320914 278695 320970 278704
rect 321098 278760 321154 278769
rect 321098 278695 321154 278704
rect 320928 269142 320956 278695
rect 320916 269136 320968 269142
rect 320914 269104 320916 269113
rect 321100 269136 321152 269142
rect 320968 269104 320970 269113
rect 320914 269039 320970 269048
rect 321098 269104 321100 269113
rect 321152 269104 321154 269113
rect 321098 269039 321154 269048
rect 320928 259486 320956 269039
rect 320916 259480 320968 259486
rect 320914 259448 320916 259457
rect 321100 259480 321152 259486
rect 320968 259448 320970 259457
rect 320914 259383 320970 259392
rect 321098 259448 321100 259457
rect 321152 259448 321154 259457
rect 321098 259383 321154 259392
rect 320928 249830 320956 259383
rect 320916 249824 320968 249830
rect 320914 249792 320916 249801
rect 321100 249824 321152 249830
rect 320968 249792 320970 249801
rect 320914 249727 320970 249736
rect 321098 249792 321100 249801
rect 321152 249792 321154 249801
rect 321098 249727 321154 249736
rect 320928 240174 320956 249727
rect 320916 240168 320968 240174
rect 320914 240136 320916 240145
rect 321100 240168 321152 240174
rect 320968 240136 320970 240145
rect 320914 240071 320970 240080
rect 321098 240136 321100 240145
rect 321152 240136 321154 240145
rect 321098 240071 321154 240080
rect 320928 230518 320956 240071
rect 320916 230512 320968 230518
rect 320914 230480 320916 230489
rect 321100 230512 321152 230518
rect 320968 230480 320970 230489
rect 320914 230415 320970 230424
rect 321098 230480 321100 230489
rect 321152 230480 321154 230489
rect 321098 230415 321154 230424
rect 320928 220862 320956 230415
rect 320916 220856 320968 220862
rect 320916 220798 320968 220804
rect 321100 220856 321152 220862
rect 321100 220798 321152 220804
rect 321112 219434 321140 220798
rect 321100 219428 321152 219434
rect 321100 219370 321152 219376
rect 321100 209840 321152 209846
rect 321100 209782 321152 209788
rect 321112 201657 321140 209782
rect 321098 201648 321154 201657
rect 321098 201583 321154 201592
rect 321098 201512 321154 201521
rect 321098 201447 321154 201456
rect 321112 200122 321140 201447
rect 321100 200116 321152 200122
rect 321100 200058 321152 200064
rect 321100 190528 321152 190534
rect 321100 190470 321152 190476
rect 321112 182345 321140 190470
rect 321098 182336 321154 182345
rect 321098 182271 321154 182280
rect 321098 182200 321154 182209
rect 321098 182135 321154 182144
rect 321112 180810 321140 182135
rect 321100 180804 321152 180810
rect 321100 180746 321152 180752
rect 321100 171148 321152 171154
rect 321100 171090 321152 171096
rect 321112 161430 321140 171090
rect 321100 161424 321152 161430
rect 321100 161366 321152 161372
rect 321100 151836 321152 151842
rect 321100 151778 321152 151784
rect 321112 143614 321140 151778
rect 320916 143608 320968 143614
rect 320916 143550 320968 143556
rect 321100 143608 321152 143614
rect 321100 143550 321152 143556
rect 320928 142225 320956 143550
rect 320914 142216 320970 142225
rect 320914 142151 320970 142160
rect 321006 141944 321062 141953
rect 321006 141879 321062 141888
rect 321020 132530 321048 141879
rect 321008 132524 321060 132530
rect 321008 132466 321060 132472
rect 321100 132524 321152 132530
rect 321100 132466 321152 132472
rect 321112 122942 321140 132466
rect 321100 122936 321152 122942
rect 321100 122878 321152 122884
rect 320916 122868 320968 122874
rect 320916 122810 320968 122816
rect 320928 113257 320956 122810
rect 320914 113248 320970 113257
rect 320914 113183 320970 113192
rect 321098 113248 321154 113257
rect 321098 113183 321154 113192
rect 321112 106078 321140 113183
rect 321100 106072 321152 106078
rect 321100 106014 321152 106020
rect 321204 103630 321232 326352
rect 321284 326334 321336 326340
rect 321192 103624 321244 103630
rect 321192 103566 321244 103572
rect 321296 103494 321324 326334
rect 321100 103488 321152 103494
rect 321100 103430 321152 103436
rect 321284 103488 321336 103494
rect 321284 103430 321336 103436
rect 321112 98682 321140 103430
rect 321284 103284 321336 103290
rect 321284 103226 321336 103232
rect 321112 98654 321232 98682
rect 321100 93900 321152 93906
rect 321100 93842 321152 93848
rect 321112 84318 321140 93842
rect 321100 84312 321152 84318
rect 321100 84254 321152 84260
rect 320824 82952 320876 82958
rect 320824 82894 320876 82900
rect 320836 82822 320864 82894
rect 320824 82816 320876 82822
rect 320824 82758 320876 82764
rect 321100 73228 321152 73234
rect 321100 73170 321152 73176
rect 321112 64818 321140 73170
rect 321020 64790 321140 64818
rect 321020 63510 321048 64790
rect 321008 63504 321060 63510
rect 321008 63446 321060 63452
rect 321100 45620 321152 45626
rect 321100 45562 321152 45568
rect 321112 45506 321140 45562
rect 321020 45478 321140 45506
rect 321020 40730 321048 45478
rect 321008 40724 321060 40730
rect 321008 40666 321060 40672
rect 321008 31748 321060 31754
rect 321008 31690 321060 31696
rect 321020 12073 321048 31690
rect 321006 12064 321062 12073
rect 321006 11999 321062 12008
rect 321204 8945 321232 98654
rect 321190 8936 321246 8945
rect 321190 8871 321246 8880
rect 320456 6996 320508 7002
rect 320456 6938 320508 6944
rect 320088 4820 320140 4826
rect 320088 4762 320140 4768
rect 320468 480 320496 6938
rect 321296 6905 321324 103226
rect 321282 6896 321338 6905
rect 321282 6831 321338 6840
rect 321388 5409 321416 330550
rect 321374 5400 321430 5409
rect 321374 5335 321430 5344
rect 321480 5273 321508 335378
rect 321572 330410 321600 340068
rect 321664 340054 321770 340082
rect 321848 340054 322046 340082
rect 322124 340054 322322 340082
rect 321664 330478 321692 340054
rect 321848 330546 321876 340054
rect 322020 337408 322072 337414
rect 322020 337350 322072 337356
rect 322032 337249 322060 337350
rect 322018 337240 322074 337249
rect 322018 337175 322074 337184
rect 322124 335594 322152 340054
rect 322204 337408 322256 337414
rect 322204 337350 322256 337356
rect 321940 335566 322152 335594
rect 321836 330540 321888 330546
rect 321836 330482 321888 330488
rect 321652 330472 321704 330478
rect 321940 330460 321968 335566
rect 322216 335458 322244 337350
rect 322124 335430 322244 335458
rect 322124 330528 322152 335430
rect 322492 335322 322520 340068
rect 322768 337414 322796 340068
rect 322952 340054 323058 340082
rect 322756 337408 322808 337414
rect 322756 337350 322808 337356
rect 322216 335294 322520 335322
rect 322216 330664 322244 335294
rect 322216 330636 322888 330664
rect 322664 330540 322716 330546
rect 322124 330500 322612 330528
rect 321940 330432 322428 330460
rect 321652 330414 321704 330420
rect 321560 330404 321612 330410
rect 321560 330346 321612 330352
rect 322400 316554 322428 330432
rect 322480 330404 322532 330410
rect 322480 330346 322532 330352
rect 322216 316526 322428 316554
rect 322216 299538 322244 316526
rect 322296 312724 322348 312730
rect 322296 312666 322348 312672
rect 322308 311166 322336 312666
rect 322296 311160 322348 311166
rect 322296 311102 322348 311108
rect 322204 299532 322256 299538
rect 322204 299474 322256 299480
rect 322296 299532 322348 299538
rect 322296 299474 322348 299480
rect 322308 293298 322336 299474
rect 322216 293270 322336 293298
rect 322216 289882 322244 293270
rect 322204 289876 322256 289882
rect 322204 289818 322256 289824
rect 322204 289740 322256 289746
rect 322204 289682 322256 289688
rect 322216 280242 322244 289682
rect 322216 280214 322336 280242
rect 322308 263634 322336 280214
rect 322296 263628 322348 263634
rect 322296 263570 322348 263576
rect 322296 259480 322348 259486
rect 322294 259448 322296 259457
rect 322348 259448 322350 259457
rect 322294 259383 322350 259392
rect 322202 259312 322258 259321
rect 322202 259247 322258 259256
rect 322216 258058 322244 259247
rect 322112 258052 322164 258058
rect 322112 257994 322164 258000
rect 322204 258052 322256 258058
rect 322204 257994 322256 258000
rect 322124 248441 322152 257994
rect 322110 248432 322166 248441
rect 322110 248367 322166 248376
rect 322294 248432 322350 248441
rect 322294 248367 322350 248376
rect 322308 238746 322336 248367
rect 322112 238740 322164 238746
rect 322112 238682 322164 238688
rect 322296 238740 322348 238746
rect 322296 238682 322348 238688
rect 322124 229129 322152 238682
rect 322110 229120 322166 229129
rect 322110 229055 322166 229064
rect 322294 229120 322350 229129
rect 322294 229055 322350 229064
rect 322308 224262 322336 229055
rect 322112 224256 322164 224262
rect 322112 224198 322164 224204
rect 322296 224256 322348 224262
rect 322296 224198 322348 224204
rect 322124 219473 322152 224198
rect 322110 219464 322166 219473
rect 322110 219399 322166 219408
rect 322294 219464 322350 219473
rect 322294 219399 322350 219408
rect 322308 219366 322336 219399
rect 322296 219360 322348 219366
rect 322296 219302 322348 219308
rect 322112 209840 322164 209846
rect 322112 209782 322164 209788
rect 322124 201521 322152 209782
rect 322110 201512 322166 201521
rect 322110 201447 322166 201456
rect 322294 201512 322350 201521
rect 322294 201447 322350 201456
rect 322308 200122 322336 201447
rect 322296 200116 322348 200122
rect 322296 200058 322348 200064
rect 322204 190528 322256 190534
rect 322204 190470 322256 190476
rect 322216 182186 322244 190470
rect 322216 182158 322336 182186
rect 322308 171222 322336 182158
rect 322296 171216 322348 171222
rect 322296 171158 322348 171164
rect 322388 171148 322440 171154
rect 322388 171090 322440 171096
rect 322400 167142 322428 171090
rect 322388 167136 322440 167142
rect 322388 167078 322440 167084
rect 322296 166932 322348 166938
rect 322296 166874 322348 166880
rect 322308 161401 322336 166874
rect 322294 161392 322350 161401
rect 322294 161327 322350 161336
rect 322386 161256 322442 161265
rect 322386 161191 322442 161200
rect 322400 151774 322428 161191
rect 322296 151768 322348 151774
rect 322296 151710 322348 151716
rect 322388 151768 322440 151774
rect 322388 151710 322440 151716
rect 322308 142118 322336 151710
rect 322296 142112 322348 142118
rect 322296 142054 322348 142060
rect 322296 141976 322348 141982
rect 322296 141918 322348 141924
rect 322308 122942 322336 141918
rect 322296 122936 322348 122942
rect 322296 122878 322348 122884
rect 322388 122732 322440 122738
rect 322388 122674 322440 122680
rect 322400 104922 322428 122674
rect 322296 104916 322348 104922
rect 322296 104858 322348 104864
rect 322388 104916 322440 104922
rect 322388 104858 322440 104864
rect 322308 103494 322336 104858
rect 322296 103488 322348 103494
rect 322296 103430 322348 103436
rect 322388 93900 322440 93906
rect 322388 93842 322440 93848
rect 322400 85610 322428 93842
rect 322296 85604 322348 85610
rect 322296 85546 322348 85552
rect 322388 85604 322440 85610
rect 322388 85546 322440 85552
rect 322308 74798 322336 85546
rect 322296 74792 322348 74798
rect 322296 74734 322348 74740
rect 322296 74656 322348 74662
rect 322296 74598 322348 74604
rect 322308 74526 322336 74598
rect 322296 74520 322348 74526
rect 322296 74462 322348 74468
rect 322388 74452 322440 74458
rect 322388 74394 322440 74400
rect 322400 64870 322428 74394
rect 322388 64864 322440 64870
rect 322388 64806 322440 64812
rect 322296 55344 322348 55350
rect 322296 55286 322348 55292
rect 322308 55214 322336 55286
rect 322296 55208 322348 55214
rect 322296 55150 322348 55156
rect 322388 55208 322440 55214
rect 322388 55150 322440 55156
rect 322400 45558 322428 55150
rect 322388 45552 322440 45558
rect 322388 45494 322440 45500
rect 322296 40724 322348 40730
rect 322296 40666 322348 40672
rect 322308 11937 322336 40666
rect 322294 11928 322350 11937
rect 322294 11863 322350 11872
rect 322492 11257 322520 330346
rect 322584 312730 322612 330500
rect 322664 330482 322716 330488
rect 322572 312724 322624 312730
rect 322572 312666 322624 312672
rect 322572 311160 322624 311166
rect 322572 311102 322624 311108
rect 322478 11248 322534 11257
rect 322478 11183 322534 11192
rect 322480 11076 322532 11082
rect 322480 11018 322532 11024
rect 321652 8968 321704 8974
rect 321652 8910 321704 8916
rect 321466 5264 321522 5273
rect 321466 5199 321522 5208
rect 321664 480 321692 8910
rect 322492 7002 322520 11018
rect 322584 8974 322612 311102
rect 322676 11082 322704 330482
rect 322756 330472 322808 330478
rect 322756 330414 322808 330420
rect 322664 11076 322716 11082
rect 322664 11018 322716 11024
rect 322768 9194 322796 330414
rect 322676 9166 322796 9194
rect 322572 8968 322624 8974
rect 322572 8910 322624 8916
rect 322480 6996 322532 7002
rect 322480 6938 322532 6944
rect 322676 5137 322704 9166
rect 322662 5128 322718 5137
rect 322662 5063 322718 5072
rect 322860 5001 322888 330636
rect 322952 330478 322980 340054
rect 323124 337476 323176 337482
rect 323124 337418 323176 337424
rect 323136 330546 323164 337418
rect 323228 330614 323256 340068
rect 323308 335028 323360 335034
rect 323308 334970 323360 334976
rect 323216 330608 323268 330614
rect 323216 330550 323268 330556
rect 323124 330540 323176 330546
rect 323124 330482 323176 330488
rect 322940 330472 322992 330478
rect 322940 330414 322992 330420
rect 322940 18080 322992 18086
rect 322940 18022 322992 18028
rect 322952 16833 322980 18022
rect 322938 16824 322994 16833
rect 322938 16759 322994 16768
rect 323320 11801 323348 334970
rect 323400 331764 323452 331770
rect 323400 331706 323452 331712
rect 323306 11792 323362 11801
rect 323306 11727 323362 11736
rect 323412 11665 323440 331706
rect 323504 330664 323532 340068
rect 323780 337482 323808 340068
rect 323872 340054 323978 340082
rect 324056 340054 324254 340082
rect 324424 340054 324530 340082
rect 324608 340054 324714 340082
rect 324884 340054 324990 340082
rect 325068 340054 325266 340082
rect 325344 340054 325450 340082
rect 325726 340054 325924 340082
rect 323768 337476 323820 337482
rect 323768 337418 323820 337424
rect 323872 331770 323900 340054
rect 323952 337476 324004 337482
rect 323952 337418 324004 337424
rect 323964 337249 323992 337418
rect 323950 337240 324006 337249
rect 323950 337175 324006 337184
rect 324056 335034 324084 340054
rect 324320 335708 324372 335714
rect 324320 335650 324372 335656
rect 324044 335028 324096 335034
rect 324044 334970 324096 334976
rect 323860 331764 323912 331770
rect 323860 331706 323912 331712
rect 323504 330636 324176 330664
rect 324044 330540 324096 330546
rect 324044 330482 324096 330488
rect 323952 330472 324004 330478
rect 323952 330414 324004 330420
rect 323964 11801 323992 330414
rect 323950 11792 324006 11801
rect 323950 11727 324006 11736
rect 324056 11665 324084 330482
rect 323398 11656 323454 11665
rect 323398 11591 323454 11600
rect 324042 11656 324098 11665
rect 324042 11591 324098 11600
rect 324044 9104 324096 9110
rect 324044 9046 324096 9052
rect 322846 4992 322902 5001
rect 322846 4927 322902 4936
rect 322846 4856 322902 4865
rect 322846 4791 322902 4800
rect 322860 480 322888 4791
rect 324056 480 324084 9046
rect 324148 8974 324176 330636
rect 324228 330608 324280 330614
rect 324228 330550 324280 330556
rect 324136 8968 324188 8974
rect 324136 8910 324188 8916
rect 324240 4865 324268 330550
rect 324226 4856 324282 4865
rect 324226 4791 324282 4800
rect 324332 3369 324360 335650
rect 324424 13025 324452 340054
rect 324608 15881 324636 340054
rect 324780 335640 324832 335646
rect 324780 335582 324832 335588
rect 324594 15872 324650 15881
rect 324594 15807 324650 15816
rect 324792 14521 324820 335582
rect 324884 18630 324912 340054
rect 325068 335714 325096 340054
rect 325056 335708 325108 335714
rect 325056 335650 325108 335656
rect 325344 335646 325372 340054
rect 325792 335708 325844 335714
rect 325792 335650 325844 335656
rect 325332 335640 325384 335646
rect 325332 335582 325384 335588
rect 324872 18624 324924 18630
rect 324872 18566 324924 18572
rect 325804 14657 325832 335650
rect 325896 335646 325924 340054
rect 325988 337385 326016 340068
rect 326172 337521 326200 340068
rect 326264 340054 326462 340082
rect 326540 340054 326738 340082
rect 326816 340054 326922 340082
rect 327198 340054 327396 340082
rect 326158 337512 326214 337521
rect 326158 337447 326214 337456
rect 325974 337376 326030 337385
rect 325974 337311 326030 337320
rect 326264 335714 326292 340054
rect 326252 335708 326304 335714
rect 326252 335650 326304 335656
rect 325884 335640 325936 335646
rect 325884 335582 325936 335588
rect 326344 335640 326396 335646
rect 326344 335582 326396 335588
rect 326356 335322 326384 335582
rect 326264 335294 326384 335322
rect 325884 335232 325936 335238
rect 325884 335174 325936 335180
rect 325896 16153 325924 335174
rect 326068 332308 326120 332314
rect 326068 332250 326120 332256
rect 325882 16144 325938 16153
rect 325882 16079 325938 16088
rect 325790 14648 325846 14657
rect 325790 14583 325846 14592
rect 324778 14512 324834 14521
rect 324778 14447 324834 14456
rect 324410 13016 324466 13025
rect 324410 12951 324466 12960
rect 324412 11144 324464 11150
rect 324412 11086 324464 11092
rect 324318 3360 324374 3369
rect 324318 3295 324374 3304
rect 324424 610 324452 11086
rect 324870 4176 324926 4185
rect 324870 4111 324926 4120
rect 324884 3738 324912 4111
rect 324872 3732 324924 3738
rect 324872 3674 324924 3680
rect 326080 3505 326108 332250
rect 326264 328506 326292 335294
rect 326540 335238 326568 340054
rect 326528 335232 326580 335238
rect 326528 335174 326580 335180
rect 326816 332314 326844 340054
rect 327264 335640 327316 335646
rect 327264 335582 327316 335588
rect 326804 332308 326856 332314
rect 326804 332250 326856 332256
rect 326252 328500 326304 328506
rect 326252 328442 326304 328448
rect 326344 328432 326396 328438
rect 326344 328374 326396 328380
rect 326356 309126 326384 328374
rect 326252 309120 326304 309126
rect 326252 309062 326304 309068
rect 326344 309120 326396 309126
rect 326344 309062 326396 309068
rect 326264 296721 326292 309062
rect 326250 296712 326306 296721
rect 326250 296647 326306 296656
rect 326434 296712 326490 296721
rect 326434 296647 326490 296656
rect 326448 287094 326476 296647
rect 326252 287088 326304 287094
rect 326252 287030 326304 287036
rect 326436 287088 326488 287094
rect 326436 287030 326488 287036
rect 326264 277409 326292 287030
rect 326250 277400 326306 277409
rect 326250 277335 326306 277344
rect 326526 277400 326582 277409
rect 326526 277335 326582 277344
rect 326540 267782 326568 277335
rect 326344 267776 326396 267782
rect 326344 267718 326396 267724
rect 326528 267776 326580 267782
rect 326528 267718 326580 267724
rect 326356 264330 326384 267718
rect 326264 264302 326384 264330
rect 326264 259434 326292 264302
rect 326264 259406 326384 259434
rect 326356 254114 326384 259406
rect 326344 254108 326396 254114
rect 326344 254050 326396 254056
rect 326252 249824 326304 249830
rect 326252 249766 326304 249772
rect 326264 230518 326292 249766
rect 326252 230512 326304 230518
rect 326252 230454 326304 230460
rect 326344 230512 326396 230518
rect 326344 230454 326396 230460
rect 326356 220930 326384 230454
rect 326344 220924 326396 220930
rect 326344 220866 326396 220872
rect 326252 220856 326304 220862
rect 326252 220798 326304 220804
rect 326264 215422 326292 220798
rect 326252 215416 326304 215422
rect 326252 215358 326304 215364
rect 326252 200184 326304 200190
rect 326252 200126 326304 200132
rect 326264 196110 326292 200126
rect 326252 196104 326304 196110
rect 326252 196046 326304 196052
rect 326252 195968 326304 195974
rect 326252 195910 326304 195916
rect 326264 174570 326292 195910
rect 326264 174542 326384 174570
rect 326356 169726 326384 174542
rect 326344 169720 326396 169726
rect 326344 169662 326396 169668
rect 326436 161356 326488 161362
rect 326436 161298 326488 161304
rect 326448 151858 326476 161298
rect 326356 151830 326476 151858
rect 326356 142186 326384 151830
rect 326160 142180 326212 142186
rect 326160 142122 326212 142128
rect 326344 142180 326396 142186
rect 326344 142122 326396 142128
rect 326172 132530 326200 142122
rect 326160 132524 326212 132530
rect 326160 132466 326212 132472
rect 326252 132524 326304 132530
rect 326252 132466 326304 132472
rect 326264 124234 326292 132466
rect 326252 124228 326304 124234
rect 326252 124170 326304 124176
rect 326344 124228 326396 124234
rect 326344 124170 326396 124176
rect 326356 114510 326384 124170
rect 326160 114504 326212 114510
rect 326160 114446 326212 114452
rect 326344 114504 326396 114510
rect 326344 114446 326396 114452
rect 326172 113150 326200 114446
rect 326160 113144 326212 113150
rect 326160 113086 326212 113092
rect 326252 103556 326304 103562
rect 326252 103498 326304 103504
rect 326264 84182 326292 103498
rect 326252 84176 326304 84182
rect 326252 84118 326304 84124
rect 326344 84176 326396 84182
rect 326344 84118 326396 84124
rect 326356 68354 326384 84118
rect 326264 68326 326384 68354
rect 326264 63510 326292 68326
rect 326252 63504 326304 63510
rect 326252 63446 326304 63452
rect 326344 63504 326396 63510
rect 326344 63446 326396 63452
rect 326356 62098 326384 63446
rect 326264 62070 326384 62098
rect 326264 52494 326292 62070
rect 326160 52488 326212 52494
rect 326160 52430 326212 52436
rect 326252 52488 326304 52494
rect 326252 52430 326304 52436
rect 326172 44266 326200 52430
rect 326160 44260 326212 44266
rect 326160 44202 326212 44208
rect 326252 44260 326304 44266
rect 326252 44202 326304 44208
rect 326264 44130 326292 44202
rect 326252 44124 326304 44130
rect 326252 44066 326304 44072
rect 326344 27668 326396 27674
rect 326344 27610 326396 27616
rect 326356 19446 326384 27610
rect 326344 19440 326396 19446
rect 326344 19382 326396 19388
rect 326160 19372 326212 19378
rect 326160 19314 326212 19320
rect 326172 16017 326200 19314
rect 326158 16008 326214 16017
rect 326158 15943 326214 15952
rect 327078 6896 327134 6905
rect 327078 6831 327134 6840
rect 326436 4208 326488 4214
rect 326436 4150 326488 4156
rect 326066 3496 326122 3505
rect 326066 3431 326122 3440
rect 324412 604 324464 610
rect 324412 546 324464 552
rect 325240 604 325292 610
rect 325240 546 325292 552
rect 325252 480 325280 546
rect 326448 480 326476 4150
rect 327092 3602 327120 6831
rect 327276 3777 327304 335582
rect 327368 335510 327396 340054
rect 327356 335504 327408 335510
rect 327356 335446 327408 335452
rect 327356 335368 327408 335374
rect 327356 335310 327408 335316
rect 327368 16425 327396 335310
rect 327354 16416 327410 16425
rect 327354 16351 327410 16360
rect 327460 16289 327488 340068
rect 327552 340054 327658 340082
rect 327828 340054 327934 340082
rect 327552 335646 327580 340054
rect 327540 335640 327592 335646
rect 327540 335582 327592 335588
rect 327540 335504 327592 335510
rect 327540 335446 327592 335452
rect 327446 16280 327502 16289
rect 327446 16215 327502 16224
rect 327262 3768 327318 3777
rect 327262 3703 327318 3712
rect 327552 3641 327580 335446
rect 327632 8356 327684 8362
rect 327632 8298 327684 8304
rect 327538 3632 327594 3641
rect 327080 3596 327132 3602
rect 327538 3567 327594 3576
rect 327080 3538 327132 3544
rect 327644 480 327672 8298
rect 327828 3466 327856 340054
rect 328196 337657 328224 340068
rect 328288 340054 328394 340082
rect 328670 340054 328776 340082
rect 328182 337648 328238 337657
rect 328182 337583 328238 337592
rect 328288 335374 328316 340054
rect 328552 335776 328604 335782
rect 328552 335718 328604 335724
rect 328460 335708 328512 335714
rect 328460 335650 328512 335656
rect 328276 335368 328328 335374
rect 328276 335310 328328 335316
rect 328472 8362 328500 335650
rect 328460 8356 328512 8362
rect 328460 8298 328512 8304
rect 328460 6996 328512 7002
rect 328460 6938 328512 6944
rect 328472 3466 328500 6938
rect 328564 4049 328592 335718
rect 328642 10976 328698 10985
rect 328642 10911 328698 10920
rect 328550 4040 328606 4049
rect 328550 3975 328606 3984
rect 328656 3534 328684 10911
rect 328748 3913 328776 340054
rect 328840 340054 328946 340082
rect 329024 340054 329130 340082
rect 329208 340054 329406 340082
rect 329576 340054 329682 340082
rect 329866 340054 330064 340082
rect 330142 340054 330248 340082
rect 328840 335782 328868 340054
rect 328828 335776 328880 335782
rect 328828 335718 328880 335724
rect 329024 335714 329052 340054
rect 329012 335708 329064 335714
rect 329012 335650 329064 335656
rect 329208 335594 329236 340054
rect 328840 335566 329236 335594
rect 328840 18057 328868 335566
rect 329576 331906 329604 340054
rect 329932 335640 329984 335646
rect 329932 335582 329984 335588
rect 329012 331900 329064 331906
rect 329012 331842 329064 331848
rect 329564 331900 329616 331906
rect 329564 331842 329616 331848
rect 329024 322266 329052 331842
rect 329024 322238 329144 322266
rect 329116 307834 329144 322238
rect 329012 307828 329064 307834
rect 329012 307770 329064 307776
rect 329104 307828 329156 307834
rect 329104 307770 329156 307776
rect 329024 298081 329052 307770
rect 329010 298072 329066 298081
rect 329010 298007 329066 298016
rect 329194 298072 329250 298081
rect 329194 298007 329250 298016
rect 329208 288522 329236 298007
rect 329012 288516 329064 288522
rect 329012 288458 329064 288464
rect 329196 288516 329248 288522
rect 329196 288458 329248 288464
rect 329024 288425 329052 288458
rect 329010 288416 329066 288425
rect 329010 288351 329066 288360
rect 329194 288416 329250 288425
rect 329194 288351 329250 288360
rect 329024 278798 329052 278829
rect 329208 278798 329236 288351
rect 329012 278792 329064 278798
rect 328932 278740 329012 278746
rect 328932 278734 329064 278740
rect 329196 278792 329248 278798
rect 329196 278734 329248 278740
rect 328932 278718 329052 278734
rect 328932 270638 328960 278718
rect 328920 270632 328972 270638
rect 328920 270574 328972 270580
rect 328920 270496 328972 270502
rect 328920 270438 328972 270444
rect 328932 260914 328960 270438
rect 328920 260908 328972 260914
rect 328920 260850 328972 260856
rect 329012 260908 329064 260914
rect 329012 260850 329064 260856
rect 329024 241618 329052 260850
rect 329024 241590 329144 241618
rect 329116 241346 329144 241590
rect 329024 241318 329144 241346
rect 329024 237386 329052 241318
rect 329012 237380 329064 237386
rect 329012 237322 329064 237328
rect 329196 237380 329248 237386
rect 329196 237322 329248 237328
rect 329208 227746 329236 237322
rect 329116 227718 329236 227746
rect 329116 216730 329144 227718
rect 329024 216702 329144 216730
rect 329024 215286 329052 216702
rect 329012 215280 329064 215286
rect 329012 215222 329064 215228
rect 329104 205692 329156 205698
rect 329104 205634 329156 205640
rect 329116 197334 329144 205634
rect 329104 197328 329156 197334
rect 329104 197270 329156 197276
rect 329012 187740 329064 187746
rect 329012 187682 329064 187688
rect 329024 179382 329052 187682
rect 329012 179376 329064 179382
rect 329012 179318 329064 179324
rect 329104 179376 329156 179382
rect 329104 179318 329156 179324
rect 329116 161498 329144 179318
rect 329012 161492 329064 161498
rect 329012 161434 329064 161440
rect 329104 161492 329156 161498
rect 329104 161434 329156 161440
rect 329024 140758 329052 161434
rect 329012 140752 329064 140758
rect 329012 140694 329064 140700
rect 329196 131164 329248 131170
rect 329196 131106 329248 131112
rect 329208 124234 329236 131106
rect 329104 124228 329156 124234
rect 329104 124170 329156 124176
rect 329196 124228 329248 124234
rect 329196 124170 329248 124176
rect 329116 114578 329144 124170
rect 329012 114572 329064 114578
rect 329012 114514 329064 114520
rect 329104 114572 329156 114578
rect 329104 114514 329156 114520
rect 329024 103630 329052 114514
rect 329012 103624 329064 103630
rect 329012 103566 329064 103572
rect 328920 103556 328972 103562
rect 328920 103498 328972 103504
rect 328932 102134 328960 103498
rect 328920 102128 328972 102134
rect 328920 102070 328972 102076
rect 329196 92540 329248 92546
rect 329196 92482 329248 92488
rect 329208 82822 329236 92482
rect 329196 82816 329248 82822
rect 329196 82758 329248 82764
rect 329012 71800 329064 71806
rect 329012 71742 329064 71748
rect 329024 62121 329052 71742
rect 329010 62112 329066 62121
rect 329010 62047 329066 62056
rect 329194 62112 329250 62121
rect 329194 62047 329250 62056
rect 329208 52494 329236 62047
rect 329012 52488 329064 52494
rect 329012 52430 329064 52436
rect 329196 52488 329248 52494
rect 329196 52430 329248 52436
rect 329024 44198 329052 52430
rect 329012 44192 329064 44198
rect 329012 44134 329064 44140
rect 329104 44192 329156 44198
rect 329104 44134 329156 44140
rect 329116 39250 329144 44134
rect 329116 39222 329236 39250
rect 329208 34513 329236 39222
rect 329194 34504 329250 34513
rect 329194 34439 329250 34448
rect 329378 34504 329434 34513
rect 329378 34439 329434 34448
rect 329208 24886 329236 24917
rect 329392 24886 329420 34439
rect 329196 24880 329248 24886
rect 329116 24828 329196 24834
rect 329116 24822 329248 24828
rect 329380 24880 329432 24886
rect 329380 24822 329432 24828
rect 329116 24806 329236 24822
rect 328826 18048 328882 18057
rect 329116 18018 329144 24806
rect 328826 17983 328882 17992
rect 329104 18012 329156 18018
rect 329104 17954 329156 17960
rect 329104 15224 329156 15230
rect 329104 15166 329156 15172
rect 328828 11212 328880 11218
rect 328828 11154 328880 11160
rect 328734 3904 328790 3913
rect 328734 3839 328790 3848
rect 328644 3528 328696 3534
rect 328644 3470 328696 3476
rect 327816 3460 327868 3466
rect 327816 3402 327868 3408
rect 328460 3460 328512 3466
rect 328460 3402 328512 3408
rect 328840 480 328868 11154
rect 328920 8356 328972 8362
rect 328920 8298 328972 8304
rect 328932 3738 328960 8298
rect 329116 6934 329144 15166
rect 329104 6928 329156 6934
rect 329104 6870 329156 6876
rect 329196 6928 329248 6934
rect 329196 6870 329248 6876
rect 328920 3732 328972 3738
rect 328920 3674 328972 3680
rect 329208 3398 329236 6870
rect 329944 3806 329972 335582
rect 330036 4214 330064 340054
rect 330116 16652 330168 16658
rect 330116 16594 330168 16600
rect 330024 4208 330076 4214
rect 330024 4150 330076 4156
rect 329932 3800 329984 3806
rect 329932 3742 329984 3748
rect 329196 3392 329248 3398
rect 329196 3334 329248 3340
rect 330128 1578 330156 16594
rect 330220 15910 330248 340054
rect 330312 340054 330418 340082
rect 330496 340054 330602 340082
rect 330772 340054 330878 340082
rect 330956 340054 331154 340082
rect 330208 15904 330260 15910
rect 330208 15846 330260 15852
rect 330312 4185 330340 340054
rect 330496 335646 330524 340054
rect 330484 335640 330536 335646
rect 330484 335582 330536 335588
rect 330772 335345 330800 340054
rect 330956 337550 330984 340054
rect 331324 337793 331352 340068
rect 331508 340054 331614 340082
rect 331692 340054 331890 340082
rect 331310 337784 331366 337793
rect 331310 337719 331366 337728
rect 330944 337544 330996 337550
rect 330944 337486 330996 337492
rect 331404 335640 331456 335646
rect 331404 335582 331456 335588
rect 330758 335336 330814 335345
rect 330758 335271 330814 335280
rect 330942 335336 330998 335345
rect 330942 335271 330998 335280
rect 330956 325718 330984 335271
rect 330760 325712 330812 325718
rect 330760 325654 330812 325660
rect 330944 325712 330996 325718
rect 330944 325654 330996 325660
rect 330772 316062 330800 325654
rect 330576 316056 330628 316062
rect 330576 315998 330628 316004
rect 330760 316056 330812 316062
rect 330760 315998 330812 316004
rect 330588 288522 330616 315998
rect 330576 288516 330628 288522
rect 330576 288458 330628 288464
rect 330484 288448 330536 288454
rect 330484 288390 330536 288396
rect 330496 280158 330524 288390
rect 330484 280152 330536 280158
rect 330484 280094 330536 280100
rect 330576 280152 330628 280158
rect 330576 280094 330628 280100
rect 330588 273986 330616 280094
rect 330496 273958 330616 273986
rect 330496 260846 330524 273958
rect 330484 260840 330536 260846
rect 330484 260782 330536 260788
rect 330576 260840 330628 260846
rect 330576 260782 330628 260788
rect 330588 247353 330616 260782
rect 330574 247344 330630 247353
rect 330574 247279 330630 247288
rect 330574 247072 330630 247081
rect 330484 247036 330536 247042
rect 330574 247007 330576 247016
rect 330484 246978 330536 246984
rect 330628 247007 330630 247016
rect 330576 246978 330628 246984
rect 330496 237386 330524 246978
rect 330392 237380 330444 237386
rect 330392 237322 330444 237328
rect 330484 237380 330536 237386
rect 330484 237322 330536 237328
rect 330404 235958 330432 237322
rect 330392 235952 330444 235958
rect 330392 235894 330444 235900
rect 330760 230104 330812 230110
rect 330760 230046 330812 230052
rect 330772 224942 330800 230046
rect 330760 224936 330812 224942
rect 330760 224878 330812 224884
rect 330944 224936 330996 224942
rect 330944 224878 330996 224884
rect 330956 215393 330984 224878
rect 330758 215384 330814 215393
rect 330758 215319 330814 215328
rect 330942 215384 330998 215393
rect 330942 215319 330998 215328
rect 330772 215286 330800 215319
rect 330760 215280 330812 215286
rect 330760 215222 330812 215228
rect 330944 215280 330996 215286
rect 330944 215222 330996 215228
rect 330956 205737 330984 215222
rect 330758 205728 330814 205737
rect 330758 205663 330814 205672
rect 330942 205728 330998 205737
rect 330942 205663 330998 205672
rect 330772 205630 330800 205663
rect 330760 205624 330812 205630
rect 330760 205566 330812 205572
rect 330576 187740 330628 187746
rect 330576 187682 330628 187688
rect 330588 180826 330616 187682
rect 330496 180798 330616 180826
rect 330496 176474 330524 180798
rect 330496 176446 330616 176474
rect 330588 160138 330616 176446
rect 330484 160132 330536 160138
rect 330484 160074 330536 160080
rect 330576 160132 330628 160138
rect 330576 160074 330628 160080
rect 330496 150414 330524 160074
rect 330484 150408 330536 150414
rect 330484 150350 330536 150356
rect 330392 140820 330444 140826
rect 330392 140762 330444 140768
rect 330404 132530 330432 140762
rect 330392 132524 330444 132530
rect 330392 132466 330444 132472
rect 330484 132524 330536 132530
rect 330484 132466 330536 132472
rect 330496 103630 330524 132466
rect 330484 103624 330536 103630
rect 330484 103566 330536 103572
rect 330392 103556 330444 103562
rect 330392 103498 330444 103504
rect 330404 93906 330432 103498
rect 330392 93900 330444 93906
rect 330392 93842 330444 93848
rect 330484 93900 330536 93906
rect 330484 93842 330536 93848
rect 330496 79234 330524 93842
rect 330496 79206 330616 79234
rect 330588 78962 330616 79206
rect 330404 78934 330616 78962
rect 330404 66298 330432 78934
rect 330392 66292 330444 66298
rect 330392 66234 330444 66240
rect 330484 66292 330536 66298
rect 330484 66234 330536 66240
rect 330496 28778 330524 66234
rect 330496 28750 330616 28778
rect 330588 16658 330616 28750
rect 331312 16720 331364 16726
rect 331312 16662 331364 16668
rect 330392 16652 330444 16658
rect 330392 16594 330444 16600
rect 330576 16652 330628 16658
rect 330576 16594 330628 16600
rect 330404 15978 330432 16594
rect 330392 15972 330444 15978
rect 330392 15914 330444 15920
rect 331324 12322 331352 16662
rect 331416 16114 331444 335582
rect 331404 16108 331456 16114
rect 331404 16050 331456 16056
rect 331508 16046 331536 340054
rect 331588 266348 331640 266354
rect 331588 266290 331640 266296
rect 331600 256737 331628 266290
rect 331586 256728 331642 256737
rect 331586 256663 331642 256672
rect 331496 16040 331548 16046
rect 331496 15982 331548 15988
rect 331324 12294 331536 12322
rect 331220 8424 331272 8430
rect 331220 8366 331272 8372
rect 330298 4176 330354 4185
rect 330298 4111 330354 4120
rect 330036 1550 330156 1578
rect 330036 480 330064 1550
rect 331232 480 331260 8366
rect 331508 7002 331536 12294
rect 331496 6996 331548 7002
rect 331496 6938 331548 6944
rect 331692 3874 331720 340054
rect 332060 331922 332088 340068
rect 332152 340054 332350 340082
rect 332152 335646 332180 340054
rect 332612 337414 332640 340068
rect 332796 337550 332824 340068
rect 332888 340054 333086 340082
rect 333256 340054 333362 340082
rect 333440 340054 333546 340082
rect 333716 340054 333822 340082
rect 332784 337544 332836 337550
rect 332784 337486 332836 337492
rect 332600 337408 332652 337414
rect 332600 337350 332652 337356
rect 332140 335640 332192 335646
rect 332140 335582 332192 335588
rect 332692 335640 332744 335646
rect 332692 335582 332744 335588
rect 331876 331894 332088 331922
rect 331876 317422 331904 331894
rect 331772 317416 331824 317422
rect 331772 317358 331824 317364
rect 331864 317416 331916 317422
rect 331864 317358 331916 317364
rect 331784 299470 331812 317358
rect 331772 299464 331824 299470
rect 331772 299406 331824 299412
rect 331864 299464 331916 299470
rect 331864 299406 331916 299412
rect 331876 289882 331904 299406
rect 331864 289876 331916 289882
rect 331864 289818 331916 289824
rect 331772 289808 331824 289814
rect 331772 289750 331824 289756
rect 331784 280158 331812 289750
rect 331772 280152 331824 280158
rect 331772 280094 331824 280100
rect 331864 280152 331916 280158
rect 331864 280094 331916 280100
rect 331876 266354 331904 280094
rect 331864 266348 331916 266354
rect 331864 266290 331916 266296
rect 331770 256728 331826 256737
rect 331770 256663 331826 256672
rect 331784 247042 331812 256663
rect 331772 247036 331824 247042
rect 331772 246978 331824 246984
rect 331956 247036 332008 247042
rect 331956 246978 332008 246984
rect 331968 237425 331996 246978
rect 331770 237416 331826 237425
rect 331770 237351 331826 237360
rect 331954 237416 332010 237425
rect 331954 237351 332010 237360
rect 331784 231878 331812 237351
rect 331772 231872 331824 231878
rect 331772 231814 331824 231820
rect 331864 231804 331916 231810
rect 331864 231746 331916 231752
rect 331876 222222 331904 231746
rect 331772 222216 331824 222222
rect 331772 222158 331824 222164
rect 331864 222216 331916 222222
rect 331864 222158 331916 222164
rect 331784 208486 331812 222158
rect 331772 208480 331824 208486
rect 331772 208422 331824 208428
rect 331864 208412 331916 208418
rect 331864 208354 331916 208360
rect 331876 197334 331904 208354
rect 331864 197328 331916 197334
rect 331864 197270 331916 197276
rect 332048 197328 332100 197334
rect 332048 197270 332100 197276
rect 332060 178090 332088 197270
rect 331864 178084 331916 178090
rect 331864 178026 331916 178032
rect 332048 178084 332100 178090
rect 332048 178026 332100 178032
rect 331876 169862 331904 178026
rect 331864 169856 331916 169862
rect 331864 169798 331916 169804
rect 331772 168428 331824 168434
rect 331772 168370 331824 168376
rect 331784 151774 331812 168370
rect 331772 151768 331824 151774
rect 331772 151710 331824 151716
rect 331772 142180 331824 142186
rect 331772 142122 331824 142128
rect 331784 140758 331812 142122
rect 331772 140752 331824 140758
rect 331772 140694 331824 140700
rect 331772 131164 331824 131170
rect 331772 131106 331824 131112
rect 331784 121446 331812 131106
rect 331772 121440 331824 121446
rect 331772 121382 331824 121388
rect 331772 111852 331824 111858
rect 331772 111794 331824 111800
rect 331784 103494 331812 111794
rect 331772 103488 331824 103494
rect 331772 103430 331824 103436
rect 331864 103488 331916 103494
rect 331864 103430 331916 103436
rect 331876 85610 331904 103430
rect 331772 85604 331824 85610
rect 331772 85546 331824 85552
rect 331864 85604 331916 85610
rect 331864 85546 331916 85552
rect 331784 75954 331812 85546
rect 331772 75948 331824 75954
rect 331772 75890 331824 75896
rect 331864 75880 331916 75886
rect 331864 75822 331916 75828
rect 331876 66298 331904 75822
rect 331772 66292 331824 66298
rect 331772 66234 331824 66240
rect 331864 66292 331916 66298
rect 331864 66234 331916 66240
rect 331784 63510 331812 66234
rect 331772 63504 331824 63510
rect 331772 63446 331824 63452
rect 331772 53848 331824 53854
rect 331772 53790 331824 53796
rect 331784 44130 331812 53790
rect 331772 44124 331824 44130
rect 331772 44066 331824 44072
rect 331956 44124 332008 44130
rect 331956 44066 332008 44072
rect 331968 16658 331996 44066
rect 332508 18080 332560 18086
rect 332508 18022 332560 18028
rect 332520 16969 332548 18022
rect 332506 16960 332562 16969
rect 332506 16895 332562 16904
rect 331864 16652 331916 16658
rect 331864 16594 331916 16600
rect 331956 16652 332008 16658
rect 331956 16594 332008 16600
rect 331876 3942 331904 16594
rect 332416 6996 332468 7002
rect 332416 6938 332468 6944
rect 331864 3936 331916 3942
rect 331864 3878 331916 3884
rect 331680 3868 331732 3874
rect 331680 3810 331732 3816
rect 332428 480 332456 6938
rect 332704 4078 332732 335582
rect 332784 16788 332836 16794
rect 332784 16730 332836 16736
rect 332796 16028 332824 16730
rect 332888 16182 332916 340054
rect 333256 334694 333284 340054
rect 333440 335646 333468 340054
rect 333428 335640 333480 335646
rect 333428 335582 333480 335588
rect 333060 334688 333112 334694
rect 333060 334630 333112 334636
rect 333244 334688 333296 334694
rect 333244 334630 333296 334636
rect 333072 317422 333100 334630
rect 333716 331906 333744 340054
rect 333244 331900 333296 331906
rect 333244 331842 333296 331848
rect 333704 331900 333756 331906
rect 333704 331842 333756 331848
rect 333256 322266 333284 331842
rect 333256 322238 333376 322266
rect 333348 317422 333376 322238
rect 333060 317416 333112 317422
rect 333060 317358 333112 317364
rect 333152 317416 333204 317422
rect 333152 317358 333204 317364
rect 333244 317416 333296 317422
rect 333244 317358 333296 317364
rect 333336 317416 333388 317422
rect 333336 317358 333388 317364
rect 333164 290018 333192 317358
rect 333256 299470 333284 317358
rect 333244 299464 333296 299470
rect 333244 299406 333296 299412
rect 333336 299464 333388 299470
rect 333336 299406 333388 299412
rect 333348 298110 333376 299406
rect 333244 298104 333296 298110
rect 333244 298046 333296 298052
rect 333336 298104 333388 298110
rect 333336 298046 333388 298052
rect 333152 290012 333204 290018
rect 333152 289954 333204 289960
rect 333152 288448 333204 288454
rect 333152 288390 333204 288396
rect 333164 273290 333192 288390
rect 333256 280158 333284 298046
rect 333244 280152 333296 280158
rect 333244 280094 333296 280100
rect 333336 280152 333388 280158
rect 333336 280094 333388 280100
rect 333152 273284 333204 273290
rect 333152 273226 333204 273232
rect 333060 273216 333112 273222
rect 333060 273158 333112 273164
rect 333072 263634 333100 273158
rect 333060 263628 333112 263634
rect 333060 263570 333112 263576
rect 333152 263560 333204 263566
rect 333152 263502 333204 263508
rect 333164 253978 333192 263502
rect 333348 260914 333376 280094
rect 333244 260908 333296 260914
rect 333244 260850 333296 260856
rect 333336 260908 333388 260914
rect 333336 260850 333388 260856
rect 333152 253972 333204 253978
rect 333152 253914 333204 253920
rect 333060 253904 333112 253910
rect 333060 253846 333112 253852
rect 333072 244322 333100 253846
rect 333256 247217 333284 260850
rect 333242 247208 333298 247217
rect 333242 247143 333298 247152
rect 333242 247072 333298 247081
rect 333242 247007 333244 247016
rect 333296 247007 333298 247016
rect 333428 247036 333480 247042
rect 333244 246978 333296 246984
rect 333428 246978 333480 246984
rect 333060 244316 333112 244322
rect 333060 244258 333112 244264
rect 333152 244248 333204 244254
rect 333152 244190 333204 244196
rect 333164 227746 333192 244190
rect 333440 237425 333468 246978
rect 333242 237416 333298 237425
rect 333242 237351 333298 237360
rect 333426 237416 333482 237425
rect 333426 237351 333482 237360
rect 333256 231826 333284 237351
rect 333256 231798 333376 231826
rect 333072 227730 333192 227746
rect 333060 227724 333192 227730
rect 333112 227718 333192 227724
rect 333060 227666 333112 227672
rect 333072 227635 333100 227666
rect 333348 222222 333376 231798
rect 333244 222216 333296 222222
rect 333244 222158 333296 222164
rect 333336 222216 333388 222222
rect 333336 222158 333388 222164
rect 333152 218068 333204 218074
rect 333152 218010 333204 218016
rect 333164 193254 333192 218010
rect 333256 218006 333284 222158
rect 333244 218000 333296 218006
rect 333244 217942 333296 217948
rect 333336 217932 333388 217938
rect 333336 217874 333388 217880
rect 333060 193248 333112 193254
rect 333060 193190 333112 193196
rect 333152 193248 333204 193254
rect 333152 193190 333204 193196
rect 333072 191826 333100 193190
rect 333060 191820 333112 191826
rect 333060 191762 333112 191768
rect 333152 191820 333204 191826
rect 333152 191762 333204 191768
rect 333164 183938 333192 191762
rect 333348 190466 333376 217874
rect 333244 190460 333296 190466
rect 333244 190402 333296 190408
rect 333336 190460 333388 190466
rect 333336 190402 333388 190408
rect 333152 183932 333204 183938
rect 333152 183874 333204 183880
rect 333152 182096 333204 182102
rect 333152 182038 333204 182044
rect 333164 76022 333192 182038
rect 333256 173942 333284 190402
rect 333244 173936 333296 173942
rect 333244 173878 333296 173884
rect 333336 173800 333388 173806
rect 333336 173742 333388 173748
rect 333348 151842 333376 173742
rect 333244 151836 333296 151842
rect 333244 151778 333296 151784
rect 333336 151836 333388 151842
rect 333336 151778 333388 151784
rect 333256 103494 333284 151778
rect 333244 103488 333296 103494
rect 333244 103430 333296 103436
rect 333336 103488 333388 103494
rect 333336 103430 333388 103436
rect 333348 85610 333376 103430
rect 333244 85604 333296 85610
rect 333244 85546 333296 85552
rect 333336 85604 333388 85610
rect 333336 85546 333388 85552
rect 333152 76016 333204 76022
rect 333152 75958 333204 75964
rect 333256 75954 333284 85546
rect 333244 75948 333296 75954
rect 333244 75890 333296 75896
rect 333152 75880 333204 75886
rect 333152 75822 333204 75828
rect 333336 75880 333388 75886
rect 333336 75822 333388 75828
rect 333164 61418 333192 75822
rect 333348 66298 333376 75822
rect 333244 66292 333296 66298
rect 333244 66234 333296 66240
rect 333336 66292 333388 66298
rect 333336 66234 333388 66240
rect 333072 61390 333192 61418
rect 333072 51134 333100 61390
rect 333060 51128 333112 51134
rect 333060 51070 333112 51076
rect 333152 50992 333204 50998
rect 333152 50934 333204 50940
rect 333164 43466 333192 50934
rect 333072 43438 333192 43466
rect 333072 29034 333100 43438
rect 333060 29028 333112 29034
rect 333060 28970 333112 28976
rect 333152 28892 333204 28898
rect 333152 28834 333204 28840
rect 332876 16176 332928 16182
rect 332876 16118 332928 16124
rect 332796 16000 332916 16028
rect 332692 4072 332744 4078
rect 332692 4014 332744 4020
rect 332888 3890 332916 16000
rect 333164 6934 333192 28834
rect 333256 14793 333284 66234
rect 333886 64016 333942 64025
rect 333886 63951 333942 63960
rect 333900 63753 333928 63951
rect 333886 63744 333942 63753
rect 333886 63679 333942 63688
rect 333886 40352 333942 40361
rect 333886 40287 333942 40296
rect 333900 40225 333928 40287
rect 333886 40216 333942 40225
rect 333886 40151 333942 40160
rect 333886 16960 333942 16969
rect 333886 16895 333942 16904
rect 333900 16697 333928 16895
rect 333886 16688 333942 16697
rect 333886 16623 333942 16632
rect 334084 16250 334112 340068
rect 334282 340054 334480 340082
rect 334164 338564 334216 338570
rect 334164 338506 334216 338512
rect 334072 16244 334124 16250
rect 334072 16186 334124 16192
rect 334176 14929 334204 338506
rect 334348 335640 334400 335646
rect 334348 335582 334400 335588
rect 334360 16318 334388 335582
rect 334348 16312 334400 16318
rect 334348 16254 334400 16260
rect 334162 14920 334218 14929
rect 334162 14855 334218 14864
rect 333242 14784 333298 14793
rect 333242 14719 333298 14728
rect 332968 6928 333020 6934
rect 332968 6870 333020 6876
rect 333152 6928 333204 6934
rect 333152 6870 333204 6876
rect 332980 4010 333008 6870
rect 334452 4146 334480 340054
rect 334544 338570 334572 340068
rect 334636 340054 334834 340082
rect 334532 338564 334584 338570
rect 334532 338506 334584 338512
rect 334636 335646 334664 340054
rect 335004 337482 335032 340068
rect 335188 340054 335294 340082
rect 335478 340054 335584 340082
rect 334992 337476 335044 337482
rect 334992 337418 335044 337424
rect 334624 335640 334676 335646
rect 334624 335582 334676 335588
rect 335188 327146 335216 340054
rect 334532 327140 334584 327146
rect 334532 327082 334584 327088
rect 335176 327140 335228 327146
rect 335176 327082 335228 327088
rect 334544 299470 334572 327082
rect 334532 299464 334584 299470
rect 334532 299406 334584 299412
rect 334624 299464 334676 299470
rect 334624 299406 334676 299412
rect 334636 289882 334664 299406
rect 334624 289876 334676 289882
rect 334624 289818 334676 289824
rect 334532 289808 334584 289814
rect 334532 289750 334584 289756
rect 334544 280158 334572 289750
rect 334532 280152 334584 280158
rect 334532 280094 334584 280100
rect 334624 280152 334676 280158
rect 334624 280094 334676 280100
rect 334636 260914 334664 280094
rect 334532 260908 334584 260914
rect 334532 260850 334584 260856
rect 334624 260908 334676 260914
rect 334624 260850 334676 260856
rect 334544 256698 334572 260850
rect 334532 256692 334584 256698
rect 334532 256634 334584 256640
rect 334532 251116 334584 251122
rect 334532 251058 334584 251064
rect 334544 216646 334572 251058
rect 334532 216640 334584 216646
rect 334532 216582 334584 216588
rect 334624 207052 334676 207058
rect 334624 206994 334676 207000
rect 334636 197334 334664 206994
rect 334624 197328 334676 197334
rect 334624 197270 334676 197276
rect 334624 187740 334676 187746
rect 334624 187682 334676 187688
rect 334636 180878 334664 187682
rect 334624 180872 334676 180878
rect 334624 180814 334676 180820
rect 334532 179512 334584 179518
rect 334532 179454 334584 179460
rect 334544 179382 334572 179454
rect 334532 179376 334584 179382
rect 334532 179318 334584 179324
rect 334532 171080 334584 171086
rect 334532 171022 334584 171028
rect 334544 151774 334572 171022
rect 334532 151768 334584 151774
rect 334532 151710 334584 151716
rect 334532 142180 334584 142186
rect 334532 142122 334584 142128
rect 334544 131322 334572 142122
rect 334544 131294 334664 131322
rect 334636 131186 334664 131294
rect 334544 131158 334664 131186
rect 334544 131102 334572 131158
rect 334532 131096 334584 131102
rect 334532 131038 334584 131044
rect 334532 121508 334584 121514
rect 334532 121450 334584 121456
rect 334544 111790 334572 121450
rect 334532 111784 334584 111790
rect 334532 111726 334584 111732
rect 334532 102264 334584 102270
rect 334532 102206 334584 102212
rect 334544 102134 334572 102206
rect 334532 102128 334584 102134
rect 334532 102070 334584 102076
rect 334624 92540 334676 92546
rect 334624 92482 334676 92488
rect 334636 66298 334664 92482
rect 334532 66292 334584 66298
rect 334532 66234 334584 66240
rect 334624 66292 334676 66298
rect 334624 66234 334676 66240
rect 334544 61470 334572 66234
rect 334532 61464 334584 61470
rect 334532 61406 334584 61412
rect 334532 46980 334584 46986
rect 334532 46922 334584 46928
rect 334544 15065 334572 46922
rect 335452 40316 335504 40322
rect 335452 40258 335504 40264
rect 335464 40225 335492 40258
rect 335450 40216 335506 40225
rect 335450 40151 335506 40160
rect 335360 16856 335412 16862
rect 335360 16798 335412 16804
rect 334530 15056 334586 15065
rect 334530 14991 334586 15000
rect 334716 8492 334768 8498
rect 334716 8434 334768 8440
rect 334440 4140 334492 4146
rect 334440 4082 334492 4088
rect 332968 4004 333020 4010
rect 332968 3946 333020 3952
rect 332888 3862 333652 3890
rect 333624 480 333652 3862
rect 334728 480 334756 8434
rect 335372 610 335400 16798
rect 335556 16386 335584 340054
rect 335740 337686 335768 340068
rect 335832 340054 336030 340082
rect 335728 337680 335780 337686
rect 335728 337622 335780 337628
rect 335832 335628 335860 340054
rect 335648 335600 335860 335628
rect 335544 16380 335596 16386
rect 335544 16322 335596 16328
rect 335648 15201 335676 335600
rect 336200 327214 336228 340068
rect 336476 337822 336504 340068
rect 336766 340054 336872 340082
rect 336950 340054 337148 340082
rect 336464 337816 336516 337822
rect 336464 337758 336516 337764
rect 336844 333946 336872 340054
rect 337016 335640 337068 335646
rect 337016 335582 337068 335588
rect 336832 333940 336884 333946
rect 336832 333882 336884 333888
rect 336832 333804 336884 333810
rect 336832 333746 336884 333752
rect 336188 327208 336240 327214
rect 336188 327150 336240 327156
rect 335820 327140 335872 327146
rect 335820 327082 335872 327088
rect 335832 325650 335860 327082
rect 335820 325644 335872 325650
rect 335820 325586 335872 325592
rect 336004 316056 336056 316062
rect 336004 315998 336056 316004
rect 336016 306406 336044 315998
rect 335820 306400 335872 306406
rect 336004 306400 336056 306406
rect 335872 306348 335952 306354
rect 335820 306342 335952 306348
rect 336004 306342 336056 306348
rect 335832 306326 335952 306342
rect 335924 296750 335952 306326
rect 335912 296744 335964 296750
rect 335912 296686 335964 296692
rect 336004 296744 336056 296750
rect 336004 296686 336056 296692
rect 336016 288522 336044 296686
rect 335820 288516 335872 288522
rect 335820 288458 335872 288464
rect 336004 288516 336056 288522
rect 336004 288458 336056 288464
rect 335832 288425 335860 288458
rect 335818 288416 335874 288425
rect 335818 288351 335874 288360
rect 336002 288416 336058 288425
rect 336002 288351 336058 288360
rect 335832 278798 335860 278829
rect 336016 278798 336044 288351
rect 335820 278792 335872 278798
rect 335740 278740 335820 278746
rect 335740 278734 335872 278740
rect 336004 278792 336056 278798
rect 336004 278734 336056 278740
rect 335740 278718 335860 278734
rect 335740 260914 335768 278718
rect 335728 260908 335780 260914
rect 335728 260850 335780 260856
rect 335820 260908 335872 260914
rect 335820 260850 335872 260856
rect 335832 258058 335860 260850
rect 335820 258052 335872 258058
rect 335820 257994 335872 258000
rect 335820 250980 335872 250986
rect 335820 250922 335872 250928
rect 335832 241534 335860 250922
rect 335820 241528 335872 241534
rect 335820 241470 335872 241476
rect 336004 241528 336056 241534
rect 336004 241470 336056 241476
rect 336016 238785 336044 241470
rect 335818 238776 335874 238785
rect 335818 238711 335874 238720
rect 336002 238776 336058 238785
rect 336002 238711 336058 238720
rect 335832 231878 335860 238711
rect 335820 231872 335872 231878
rect 335820 231814 335872 231820
rect 335912 231804 335964 231810
rect 335912 231746 335964 231752
rect 335924 218074 335952 231746
rect 335820 218068 335872 218074
rect 335820 218010 335872 218016
rect 335912 218068 335964 218074
rect 335912 218010 335964 218016
rect 335832 209778 335860 218010
rect 335820 209772 335872 209778
rect 335820 209714 335872 209720
rect 336096 203584 336148 203590
rect 336096 203526 336148 203532
rect 336108 190505 336136 203526
rect 335910 190496 335966 190505
rect 335832 190466 335910 190482
rect 335820 190460 335910 190466
rect 335872 190454 335910 190460
rect 335910 190431 335966 190440
rect 336094 190496 336150 190505
rect 336094 190431 336150 190440
rect 335820 190402 335872 190408
rect 335832 190371 335860 190402
rect 335820 180872 335872 180878
rect 335820 180814 335872 180820
rect 335832 173942 335860 180814
rect 335820 173936 335872 173942
rect 335820 173878 335872 173884
rect 335912 173800 335964 173806
rect 335912 173742 335964 173748
rect 335924 166326 335952 173742
rect 335912 166320 335964 166326
rect 335912 166262 335964 166268
rect 336096 166320 336148 166326
rect 336096 166262 336148 166268
rect 336108 161537 336136 166262
rect 335910 161528 335966 161537
rect 335832 161486 335910 161514
rect 335832 140758 335860 161486
rect 335910 161463 335966 161472
rect 336094 161528 336150 161537
rect 336094 161463 336150 161472
rect 335820 140752 335872 140758
rect 335820 140694 335872 140700
rect 335912 131164 335964 131170
rect 335912 131106 335964 131112
rect 335924 122942 335952 131106
rect 335728 122936 335780 122942
rect 335728 122878 335780 122884
rect 335912 122936 335964 122942
rect 335912 122878 335964 122884
rect 335740 122806 335768 122878
rect 335728 122800 335780 122806
rect 335728 122742 335780 122748
rect 335820 122800 335872 122806
rect 335820 122742 335872 122748
rect 335832 113150 335860 122742
rect 335820 113144 335872 113150
rect 335820 113086 335872 113092
rect 335820 103624 335872 103630
rect 335820 103566 335872 103572
rect 335832 103494 335860 103566
rect 335820 103488 335872 103494
rect 335820 103430 335872 103436
rect 335912 93900 335964 93906
rect 335912 93842 335964 93848
rect 335924 66298 335952 93842
rect 335820 66292 335872 66298
rect 335820 66234 335872 66240
rect 335912 66292 335964 66298
rect 335912 66234 335964 66240
rect 335832 16454 335860 66234
rect 336740 16924 336792 16930
rect 336740 16866 336792 16872
rect 335820 16448 335872 16454
rect 335820 16390 335872 16396
rect 335634 15192 335690 15201
rect 335634 15127 335690 15136
rect 336752 610 336780 16866
rect 336844 14550 336872 333746
rect 337028 16590 337056 335582
rect 337016 16584 337068 16590
rect 337016 16526 337068 16532
rect 337120 16522 337148 340054
rect 337108 16516 337160 16522
rect 337108 16458 337160 16464
rect 336832 14544 336884 14550
rect 336832 14486 336884 14492
rect 337212 3670 337240 340068
rect 337396 340054 337502 340082
rect 337580 340054 337686 340082
rect 337292 333940 337344 333946
rect 337292 333882 337344 333888
rect 337304 14482 337332 333882
rect 337396 333810 337424 340054
rect 337580 335646 337608 340054
rect 337948 337754 337976 340068
rect 337936 337748 337988 337754
rect 337936 337690 337988 337696
rect 337568 335640 337620 335646
rect 337568 335582 337620 335588
rect 337384 333804 337436 333810
rect 337384 333746 337436 333752
rect 337934 29336 337990 29345
rect 338118 29336 338174 29345
rect 337990 29294 338118 29322
rect 337934 29271 337990 29280
rect 338118 29271 338174 29280
rect 338224 14618 338252 340068
rect 338304 335708 338356 335714
rect 338304 335650 338356 335656
rect 338316 14686 338344 335650
rect 338408 17241 338436 340068
rect 338592 340054 338698 340082
rect 338776 340054 338974 340082
rect 339052 340054 339158 340082
rect 338488 335640 338540 335646
rect 338488 335582 338540 335588
rect 338500 18698 338528 335582
rect 338488 18692 338540 18698
rect 338488 18634 338540 18640
rect 338394 17232 338450 17241
rect 338394 17167 338450 17176
rect 338304 14680 338356 14686
rect 338304 14622 338356 14628
rect 338212 14612 338264 14618
rect 338212 14554 338264 14560
rect 337292 14476 337344 14482
rect 337292 14418 337344 14424
rect 338304 8560 338356 8566
rect 338304 8502 338356 8508
rect 337200 3664 337252 3670
rect 337200 3606 337252 3612
rect 335360 604 335412 610
rect 335360 546 335412 552
rect 335912 604 335964 610
rect 335912 546 335964 552
rect 336740 604 336792 610
rect 336740 546 336792 552
rect 337108 604 337160 610
rect 337108 546 337160 552
rect 335924 480 335952 546
rect 337120 480 337148 546
rect 338316 480 338344 8502
rect 338592 3330 338620 340054
rect 338776 335714 338804 340054
rect 338764 335708 338816 335714
rect 338764 335650 338816 335656
rect 339052 335646 339080 340054
rect 339420 337890 339448 340068
rect 339604 340054 339710 340082
rect 339408 337884 339460 337890
rect 339408 337826 339460 337832
rect 339500 335708 339552 335714
rect 339500 335650 339552 335656
rect 339040 335640 339092 335646
rect 339040 335582 339092 335588
rect 338580 3324 338632 3330
rect 338580 3266 338632 3272
rect 339512 3262 339540 335650
rect 339604 14754 339632 340054
rect 339776 335640 339828 335646
rect 339776 335582 339828 335588
rect 339788 18834 339816 335582
rect 339776 18828 339828 18834
rect 339776 18770 339828 18776
rect 339880 18766 339908 340068
rect 339972 340054 340170 340082
rect 340340 340054 340446 340082
rect 340524 340054 340630 340082
rect 339972 335714 340000 340054
rect 339960 335708 340012 335714
rect 339960 335650 340012 335656
rect 340340 328522 340368 340054
rect 340524 335646 340552 340054
rect 340892 337958 340920 340068
rect 341182 340054 341288 340082
rect 341064 338428 341116 338434
rect 341064 338370 341116 338376
rect 340880 337952 340932 337958
rect 340880 337894 340932 337900
rect 340512 335640 340564 335646
rect 340512 335582 340564 335588
rect 340972 335640 341024 335646
rect 340972 335582 341024 335588
rect 340156 328494 340368 328522
rect 340156 317422 340184 328494
rect 340144 317416 340196 317422
rect 340144 317358 340196 317364
rect 339960 307828 340012 307834
rect 339960 307770 340012 307776
rect 339972 302138 340000 307770
rect 339972 302110 340184 302138
rect 340156 299470 340184 302110
rect 339960 299464 340012 299470
rect 339960 299406 340012 299412
rect 340144 299464 340196 299470
rect 340144 299406 340196 299412
rect 339972 298110 340000 299406
rect 339960 298104 340012 298110
rect 339960 298046 340012 298052
rect 340052 282872 340104 282878
rect 340052 282814 340104 282820
rect 340064 280242 340092 282814
rect 340064 280214 340184 280242
rect 340156 280158 340184 280214
rect 340052 280152 340104 280158
rect 340052 280094 340104 280100
rect 340144 280152 340196 280158
rect 340144 280094 340196 280100
rect 340064 270745 340092 280094
rect 340050 270736 340106 270745
rect 340050 270671 340106 270680
rect 340326 270464 340382 270473
rect 340326 270399 340382 270408
rect 340340 253892 340368 270399
rect 340064 253864 340368 253892
rect 340064 244322 340092 253864
rect 340052 244316 340104 244322
rect 340052 244258 340104 244264
rect 340144 244180 340196 244186
rect 340144 244122 340196 244128
rect 340156 230586 340184 244122
rect 340144 230580 340196 230586
rect 340144 230522 340196 230528
rect 339960 230512 340012 230518
rect 339958 230480 339960 230489
rect 340012 230480 340014 230489
rect 339958 230415 340014 230424
rect 340142 230480 340198 230489
rect 340142 230415 340198 230424
rect 340156 229090 340184 230415
rect 340144 229084 340196 229090
rect 340144 229026 340196 229032
rect 340052 220788 340104 220794
rect 340052 220730 340104 220736
rect 340064 211138 340092 220730
rect 340052 211132 340104 211138
rect 340052 211074 340104 211080
rect 340236 204944 340288 204950
rect 340236 204886 340288 204892
rect 340248 195956 340276 204886
rect 340156 195928 340276 195956
rect 340156 186402 340184 195928
rect 340064 186374 340184 186402
rect 340064 178838 340092 186374
rect 340052 178832 340104 178838
rect 340052 178774 340104 178780
rect 340144 178764 340196 178770
rect 340144 178706 340196 178712
rect 340156 169114 340184 178706
rect 340144 169108 340196 169114
rect 340144 169050 340196 169056
rect 340328 169108 340380 169114
rect 340328 169050 340380 169056
rect 340340 164257 340368 169050
rect 340142 164248 340198 164257
rect 340052 164212 340104 164218
rect 340142 164183 340144 164192
rect 340052 164154 340104 164160
rect 340196 164183 340198 164192
rect 340326 164248 340382 164257
rect 340326 164183 340382 164192
rect 340144 164154 340196 164160
rect 340064 154714 340092 164154
rect 340064 154686 340184 154714
rect 340156 149818 340184 154686
rect 340156 149790 340460 149818
rect 340432 144945 340460 149790
rect 340142 144936 340198 144945
rect 340142 144871 340198 144880
rect 340418 144936 340474 144945
rect 340418 144871 340474 144880
rect 340156 135318 340184 144871
rect 340144 135312 340196 135318
rect 340144 135254 340196 135260
rect 340052 135244 340104 135250
rect 340052 135186 340104 135192
rect 340064 133890 340092 135186
rect 340052 133884 340104 133890
rect 340052 133826 340104 133832
rect 340144 124228 340196 124234
rect 340144 124170 340196 124176
rect 340156 115530 340184 124170
rect 340144 115524 340196 115530
rect 340144 115466 340196 115472
rect 340052 108996 340104 109002
rect 340052 108938 340104 108944
rect 340064 106298 340092 108938
rect 340064 106270 340184 106298
rect 340156 96642 340184 106270
rect 340064 96614 340184 96642
rect 340064 95198 340092 96614
rect 340052 95192 340104 95198
rect 340052 95134 340104 95140
rect 340144 85604 340196 85610
rect 340144 85546 340196 85552
rect 340156 85490 340184 85546
rect 340156 85462 340276 85490
rect 340248 75970 340276 85462
rect 340156 75942 340276 75970
rect 340156 71074 340184 75942
rect 340156 71046 340276 71074
rect 340248 51066 340276 71046
rect 340052 51060 340104 51066
rect 340052 51002 340104 51008
rect 340236 51060 340288 51066
rect 340236 51002 340288 51008
rect 340064 28966 340092 51002
rect 340052 28960 340104 28966
rect 340052 28902 340104 28908
rect 339960 28892 340012 28898
rect 339960 28834 340012 28840
rect 339868 18760 339920 18766
rect 339868 18702 339920 18708
rect 339776 17060 339828 17066
rect 339776 17002 339828 17008
rect 339684 16992 339736 16998
rect 339684 16934 339736 16940
rect 339592 14748 339644 14754
rect 339592 14690 339644 14696
rect 339696 7002 339724 16934
rect 339684 6996 339736 7002
rect 339684 6938 339736 6944
rect 339500 3256 339552 3262
rect 339500 3198 339552 3204
rect 339788 1306 339816 17002
rect 339972 14822 340000 28834
rect 340984 14958 341012 335582
rect 341076 18902 341104 338370
rect 341064 18896 341116 18902
rect 341064 18838 341116 18844
rect 340972 14952 341024 14958
rect 340972 14894 341024 14900
rect 341260 14890 341288 340054
rect 341352 338434 341380 340068
rect 341340 338428 341392 338434
rect 341340 338370 341392 338376
rect 341628 338094 341656 340068
rect 341720 340054 341918 340082
rect 341616 338088 341668 338094
rect 341616 338030 341668 338036
rect 341720 335646 341748 340054
rect 341708 335640 341760 335646
rect 341708 335582 341760 335588
rect 342088 330682 342116 340068
rect 342378 340054 342576 340082
rect 342654 340054 342760 340082
rect 342444 335640 342496 335646
rect 342444 335582 342496 335588
rect 342548 335594 342576 340054
rect 342732 335714 342760 340054
rect 342720 335708 342772 335714
rect 342720 335650 342772 335656
rect 341524 330676 341576 330682
rect 341524 330618 341576 330624
rect 342076 330676 342128 330682
rect 342076 330618 342128 330624
rect 341536 328438 341564 330618
rect 341524 328432 341576 328438
rect 341524 328374 341576 328380
rect 341708 328432 341760 328438
rect 341708 328374 341760 328380
rect 341720 327078 341748 328374
rect 341708 327072 341760 327078
rect 341708 327014 341760 327020
rect 341616 317484 341668 317490
rect 341616 317426 341668 317432
rect 341628 317370 341656 317426
rect 341536 317342 341656 317370
rect 341536 311930 341564 317342
rect 341536 311902 341656 311930
rect 341628 302258 341656 311902
rect 341616 302252 341668 302258
rect 341616 302194 341668 302200
rect 341708 302116 341760 302122
rect 341708 302058 341760 302064
rect 341720 299470 341748 302058
rect 341708 299464 341760 299470
rect 341708 299406 341760 299412
rect 341708 299328 341760 299334
rect 341708 299270 341760 299276
rect 341720 282826 341748 299270
rect 341628 282798 341748 282826
rect 341628 273358 341656 282798
rect 341616 273352 341668 273358
rect 341616 273294 341668 273300
rect 341616 273216 341668 273222
rect 341616 273158 341668 273164
rect 341628 260846 341656 273158
rect 341616 260840 341668 260846
rect 341616 260782 341668 260788
rect 341708 251252 341760 251258
rect 341708 251194 341760 251200
rect 341720 244202 341748 251194
rect 341628 244174 341748 244202
rect 341628 235362 341656 244174
rect 341628 235334 341748 235362
rect 341720 216034 341748 235334
rect 341708 216028 341760 216034
rect 341708 215970 341760 215976
rect 341892 216028 341944 216034
rect 341892 215970 341944 215976
rect 341904 211177 341932 215970
rect 341706 211168 341762 211177
rect 341706 211103 341762 211112
rect 341890 211168 341946 211177
rect 341890 211103 341946 211112
rect 341720 205578 341748 211103
rect 341628 205550 341748 205578
rect 341628 196058 341656 205550
rect 341536 196030 341656 196058
rect 341536 195974 341564 196030
rect 341524 195968 341576 195974
rect 341524 195910 341576 195916
rect 341708 195968 341760 195974
rect 341708 195910 341760 195916
rect 341720 183598 341748 195910
rect 341616 183592 341668 183598
rect 341616 183534 341668 183540
rect 341708 183592 341760 183598
rect 341708 183534 341760 183540
rect 341628 166954 341656 183534
rect 341444 166926 341656 166954
rect 341444 154578 341472 166926
rect 341444 154550 341748 154578
rect 341720 147642 341748 154550
rect 341628 147614 341748 147642
rect 341628 140026 341656 147614
rect 341628 139998 341748 140026
rect 341720 128330 341748 139998
rect 341628 128302 341748 128330
rect 341628 120714 341656 128302
rect 341628 120686 341748 120714
rect 341720 109018 341748 120686
rect 341628 108990 341748 109018
rect 341628 101402 341656 108990
rect 341628 101374 341748 101402
rect 341720 75954 341748 101374
rect 341432 75948 341484 75954
rect 341432 75890 341484 75896
rect 341708 75948 341760 75954
rect 341708 75890 341760 75896
rect 341444 70394 341472 75890
rect 341444 70366 341656 70394
rect 341628 62778 341656 70366
rect 341628 62750 341748 62778
rect 341720 46986 341748 62750
rect 341524 46980 341576 46986
rect 341524 46922 341576 46928
rect 341708 46980 341760 46986
rect 341708 46922 341760 46928
rect 341536 46866 341564 46922
rect 341536 46838 341656 46866
rect 341628 22250 341656 46838
rect 341444 22222 341656 22250
rect 341444 22114 341472 22222
rect 341352 22086 341472 22114
rect 341352 18970 341380 22086
rect 341340 18964 341392 18970
rect 341340 18906 341392 18912
rect 342456 15842 342484 335582
rect 342548 335566 342760 335594
rect 342536 335504 342588 335510
rect 342536 335446 342588 335452
rect 342548 19106 342576 335446
rect 342536 19100 342588 19106
rect 342536 19042 342588 19048
rect 342444 15836 342496 15842
rect 342444 15778 342496 15784
rect 341248 14884 341300 14890
rect 341248 14826 341300 14832
rect 339960 14816 340012 14822
rect 339960 14758 340012 14764
rect 342628 12504 342680 12510
rect 342628 12446 342680 12452
rect 341892 8628 341944 8634
rect 341892 8570 341944 8576
rect 340696 6996 340748 7002
rect 340696 6938 340748 6944
rect 339512 1278 339816 1306
rect 339512 480 339540 1278
rect 340708 480 340736 6938
rect 341904 480 341932 8570
rect 342640 3074 342668 12446
rect 342732 3194 342760 335566
rect 342824 19038 342852 340068
rect 343100 338026 343128 340068
rect 343192 340054 343390 340082
rect 343468 340054 343574 340082
rect 343850 340054 344048 340082
rect 343088 338020 343140 338026
rect 343088 337962 343140 337968
rect 342904 335708 342956 335714
rect 342904 335650 342956 335656
rect 342812 19032 342864 19038
rect 342812 18974 342864 18980
rect 342916 15026 342944 335650
rect 343192 335646 343220 340054
rect 343180 335640 343232 335646
rect 343180 335582 343232 335588
rect 343468 335510 343496 340054
rect 343732 338700 343784 338706
rect 343732 338642 343784 338648
rect 343456 335504 343508 335510
rect 343456 335446 343508 335452
rect 343744 15774 343772 338642
rect 343916 335640 343968 335646
rect 343916 335582 343968 335588
rect 343928 19174 343956 335582
rect 343916 19168 343968 19174
rect 343916 19110 343968 19116
rect 343732 15768 343784 15774
rect 343732 15710 343784 15716
rect 342904 15020 342956 15026
rect 342904 14962 342956 14968
rect 342720 3188 342772 3194
rect 342720 3130 342772 3136
rect 344020 3126 344048 340054
rect 344112 338706 344140 340068
rect 344204 340054 344310 340082
rect 344100 338700 344152 338706
rect 344100 338642 344152 338648
rect 344204 335646 344232 340054
rect 344572 337346 344600 340068
rect 344664 340054 344862 340082
rect 344560 337340 344612 337346
rect 344560 337282 344612 337288
rect 344192 335640 344244 335646
rect 344192 335582 344244 335588
rect 344664 333282 344692 340054
rect 345032 335646 345060 340068
rect 345204 335708 345256 335714
rect 345204 335650 345256 335656
rect 345020 335640 345072 335646
rect 345020 335582 345072 335588
rect 345112 335572 345164 335578
rect 345112 335514 345164 335520
rect 344296 333254 344692 333282
rect 344296 328438 344324 333254
rect 344284 328432 344336 328438
rect 344284 328374 344336 328380
rect 344376 318844 344428 318850
rect 344376 318786 344428 318792
rect 344388 311914 344416 318786
rect 344192 311908 344244 311914
rect 344192 311850 344244 311856
rect 344376 311908 344428 311914
rect 344376 311850 344428 311856
rect 344204 302274 344232 311850
rect 344112 302246 344232 302274
rect 344112 302138 344140 302246
rect 344112 302110 344232 302138
rect 344204 292618 344232 302110
rect 344204 292590 344324 292618
rect 344296 275346 344324 292590
rect 344112 275318 344324 275346
rect 344112 273170 344140 275318
rect 344112 273142 344232 273170
rect 344204 263650 344232 273142
rect 344112 263622 344232 263650
rect 344112 263514 344140 263622
rect 344112 263486 344324 263514
rect 344296 244322 344324 263486
rect 344100 244316 344152 244322
rect 344100 244258 344152 244264
rect 344284 244316 344336 244322
rect 344284 244258 344336 244264
rect 344112 244202 344140 244258
rect 344112 244174 344232 244202
rect 344204 234682 344232 244174
rect 344204 234654 344324 234682
rect 344296 225010 344324 234654
rect 344100 225004 344152 225010
rect 344100 224946 344152 224952
rect 344284 225004 344336 225010
rect 344284 224946 344336 224952
rect 344112 224890 344140 224946
rect 344112 224862 344324 224890
rect 344296 205698 344324 224862
rect 344100 205692 344152 205698
rect 344100 205634 344152 205640
rect 344284 205692 344336 205698
rect 344284 205634 344336 205640
rect 344112 205578 344140 205634
rect 344112 205550 344232 205578
rect 344204 196058 344232 205550
rect 344204 196030 344324 196058
rect 344296 176746 344324 196030
rect 344296 176718 344416 176746
rect 344388 176610 344416 176718
rect 344204 176582 344416 176610
rect 344204 167090 344232 176582
rect 344112 167062 344232 167090
rect 344112 166954 344140 167062
rect 344112 166926 344232 166954
rect 344204 159338 344232 166926
rect 344204 159310 344324 159338
rect 344296 147694 344324 159310
rect 344100 147688 344152 147694
rect 344284 147688 344336 147694
rect 344152 147636 344232 147642
rect 344100 147630 344232 147636
rect 344284 147630 344336 147636
rect 344112 147614 344232 147630
rect 344204 140026 344232 147614
rect 344204 139998 344416 140026
rect 344388 137986 344416 139998
rect 344296 137958 344416 137986
rect 344296 128382 344324 137958
rect 344100 128376 344152 128382
rect 344284 128376 344336 128382
rect 344152 128324 344232 128330
rect 344100 128318 344232 128324
rect 344284 128318 344336 128324
rect 344112 128302 344232 128318
rect 344204 120714 344232 128302
rect 344204 120686 344416 120714
rect 344388 118674 344416 120686
rect 344296 118646 344416 118674
rect 344296 109070 344324 118646
rect 344100 109064 344152 109070
rect 344284 109064 344336 109070
rect 344152 109012 344232 109018
rect 344100 109006 344232 109012
rect 344284 109006 344336 109012
rect 344112 108990 344232 109006
rect 344204 101402 344232 108990
rect 344204 101374 344324 101402
rect 344296 89758 344324 101374
rect 344100 89752 344152 89758
rect 344284 89752 344336 89758
rect 344152 89700 344232 89706
rect 344100 89694 344232 89700
rect 344284 89694 344336 89700
rect 344112 89678 344232 89694
rect 344204 89570 344232 89678
rect 344204 89542 344324 89570
rect 344296 48346 344324 89542
rect 344192 48340 344244 48346
rect 344192 48282 344244 48288
rect 344284 48340 344336 48346
rect 344284 48282 344336 48288
rect 344204 41478 344232 48282
rect 344192 41472 344244 41478
rect 344192 41414 344244 41420
rect 344100 41404 344152 41410
rect 344100 41346 344152 41352
rect 344112 33810 344140 41346
rect 344926 40352 344982 40361
rect 344926 40287 344928 40296
rect 344980 40287 344982 40296
rect 344928 40258 344980 40264
rect 344112 33782 344324 33810
rect 344296 31634 344324 33782
rect 344204 31606 344324 31634
rect 344204 19378 344232 31606
rect 344100 19372 344152 19378
rect 344100 19314 344152 19320
rect 344192 19372 344244 19378
rect 344192 19314 344244 19320
rect 344112 15706 344140 19314
rect 345018 16280 345074 16289
rect 345018 16215 345020 16224
rect 345072 16215 345074 16224
rect 345020 16186 345072 16192
rect 344100 15700 344152 15706
rect 344100 15642 344152 15648
rect 345124 15638 345152 335514
rect 345112 15632 345164 15638
rect 345112 15574 345164 15580
rect 345216 15570 345244 335650
rect 345308 333282 345336 340068
rect 345400 340054 345598 340082
rect 345400 335578 345428 340054
rect 345768 337074 345796 340068
rect 346044 337278 346072 340068
rect 346136 340054 346334 340082
rect 346518 340054 346624 340082
rect 346032 337272 346084 337278
rect 346032 337214 346084 337220
rect 345756 337068 345808 337074
rect 345756 337010 345808 337016
rect 346136 335714 346164 340054
rect 346124 335708 346176 335714
rect 346124 335650 346176 335656
rect 345664 335640 345716 335646
rect 345664 335582 345716 335588
rect 345388 335572 345440 335578
rect 345388 335514 345440 335520
rect 345308 333254 345520 333282
rect 345492 331106 345520 333254
rect 345400 331078 345520 331106
rect 345400 299470 345428 331078
rect 345388 299464 345440 299470
rect 345388 299406 345440 299412
rect 345388 299328 345440 299334
rect 345388 299270 345440 299276
rect 345400 280106 345428 299270
rect 345308 280078 345428 280106
rect 345308 270570 345336 280078
rect 345296 270564 345348 270570
rect 345296 270506 345348 270512
rect 345388 270564 345440 270570
rect 345388 270506 345440 270512
rect 345400 260846 345428 270506
rect 345388 260840 345440 260846
rect 345388 260782 345440 260788
rect 345388 260704 345440 260710
rect 345388 260646 345440 260652
rect 345400 259457 345428 260646
rect 345386 259448 345442 259457
rect 345386 259383 345442 259392
rect 345570 259448 345626 259457
rect 345570 259383 345626 259392
rect 345584 249830 345612 259383
rect 345388 249824 345440 249830
rect 345388 249766 345440 249772
rect 345572 249824 345624 249830
rect 345572 249766 345624 249772
rect 345400 201482 345428 249766
rect 345388 201476 345440 201482
rect 345388 201418 345440 201424
rect 345572 201476 345624 201482
rect 345572 201418 345624 201424
rect 345584 191865 345612 201418
rect 345386 191856 345442 191865
rect 345386 191791 345442 191800
rect 345570 191856 345626 191865
rect 345570 191791 345626 191800
rect 345400 183666 345428 191791
rect 345388 183660 345440 183666
rect 345388 183602 345440 183608
rect 345296 183592 345348 183598
rect 345296 183534 345348 183540
rect 345308 173942 345336 183534
rect 345296 173936 345348 173942
rect 345296 173878 345348 173884
rect 345388 173936 345440 173942
rect 345388 173878 345440 173884
rect 345400 164218 345428 173878
rect 345388 164212 345440 164218
rect 345388 164154 345440 164160
rect 345572 164212 345624 164218
rect 345572 164154 345624 164160
rect 345584 154601 345612 164154
rect 345386 154592 345442 154601
rect 345386 154527 345442 154536
rect 345570 154592 345626 154601
rect 345570 154527 345626 154536
rect 345400 144974 345428 154527
rect 345296 144968 345348 144974
rect 345296 144910 345348 144916
rect 345388 144968 345440 144974
rect 345388 144910 345440 144916
rect 345308 135318 345336 144910
rect 345296 135312 345348 135318
rect 345296 135254 345348 135260
rect 345388 135312 345440 135318
rect 345388 135254 345440 135260
rect 345400 133890 345428 135254
rect 345388 133884 345440 133890
rect 345388 133826 345440 133832
rect 345572 133884 345624 133890
rect 345572 133826 345624 133832
rect 345584 124273 345612 133826
rect 345294 124264 345350 124273
rect 345294 124199 345350 124208
rect 345570 124264 345626 124273
rect 345570 124199 345626 124208
rect 345308 124166 345336 124199
rect 345296 124160 345348 124166
rect 345296 124102 345348 124108
rect 345388 124092 345440 124098
rect 345388 124034 345440 124040
rect 345400 106298 345428 124034
rect 345308 106270 345428 106298
rect 345308 96694 345336 106270
rect 345296 96688 345348 96694
rect 345296 96630 345348 96636
rect 345388 96688 345440 96694
rect 345388 96630 345440 96636
rect 345400 67590 345428 96630
rect 345388 67584 345440 67590
rect 345388 67526 345440 67532
rect 345388 57996 345440 58002
rect 345388 57938 345440 57944
rect 345400 48414 345428 57938
rect 345388 48408 345440 48414
rect 345388 48350 345440 48356
rect 345296 48340 345348 48346
rect 345296 48282 345348 48288
rect 345308 38690 345336 48282
rect 345296 38684 345348 38690
rect 345296 38626 345348 38632
rect 345388 38684 345440 38690
rect 345388 38626 345440 38632
rect 345400 19378 345428 38626
rect 345388 19372 345440 19378
rect 345388 19314 345440 19320
rect 345480 19372 345532 19378
rect 345480 19314 345532 19320
rect 345492 17898 345520 19314
rect 345676 19242 345704 335582
rect 346596 19310 346624 340054
rect 346688 340054 346794 340082
rect 346964 340054 347070 340082
rect 346584 19304 346636 19310
rect 346584 19246 346636 19252
rect 345664 19236 345716 19242
rect 345664 19178 345716 19184
rect 345400 17870 345520 17898
rect 345204 15564 345256 15570
rect 345204 15506 345256 15512
rect 345400 11082 345428 17870
rect 346398 16552 346454 16561
rect 346398 16487 346454 16496
rect 346412 16250 346440 16487
rect 346400 16244 346452 16250
rect 346400 16186 346452 16192
rect 346584 12572 346636 12578
rect 346584 12514 346636 12520
rect 345388 11076 345440 11082
rect 345388 11018 345440 11024
rect 345480 8696 345532 8702
rect 345480 8638 345532 8644
rect 345388 8356 345440 8362
rect 345388 8298 345440 8304
rect 344284 5568 344336 5574
rect 344284 5510 344336 5516
rect 344008 3120 344060 3126
rect 342640 3046 343128 3074
rect 344008 3062 344060 3068
rect 343100 480 343128 3046
rect 344296 480 344324 5510
rect 345400 3058 345428 8298
rect 345388 3052 345440 3058
rect 345388 2994 345440 3000
rect 345492 480 345520 8638
rect 346596 2802 346624 12514
rect 346688 2922 346716 340054
rect 346964 15502 346992 340054
rect 347240 337006 347268 340068
rect 347516 337210 347544 340068
rect 347504 337204 347556 337210
rect 347504 337146 347556 337152
rect 347228 337000 347280 337006
rect 347228 336942 347280 336948
rect 347792 335646 347820 340068
rect 347884 340054 347990 340082
rect 347780 335640 347832 335646
rect 347780 335582 347832 335588
rect 346952 15496 347004 15502
rect 346952 15438 347004 15444
rect 347884 5794 347912 340054
rect 348056 335708 348108 335714
rect 348056 335650 348108 335656
rect 348068 15366 348096 335650
rect 348252 331242 348280 340068
rect 348344 340054 348542 340082
rect 348344 335714 348372 340054
rect 348712 336938 348740 340068
rect 348988 337142 349016 340068
rect 349278 340054 349384 340082
rect 348976 337136 349028 337142
rect 348976 337078 349028 337084
rect 348700 336932 348752 336938
rect 348700 336874 348752 336880
rect 348332 335708 348384 335714
rect 348332 335650 348384 335656
rect 348424 335640 348476 335646
rect 348424 335582 348476 335588
rect 348160 331214 348280 331242
rect 348056 15360 348108 15366
rect 348056 15302 348108 15308
rect 347792 5766 347912 5794
rect 346676 2916 346728 2922
rect 346676 2858 346728 2864
rect 347792 2854 347820 5766
rect 347872 5636 347924 5642
rect 347872 5578 347924 5584
rect 347780 2848 347832 2854
rect 346596 2774 346716 2802
rect 347780 2790 347832 2796
rect 346688 480 346716 2774
rect 347884 480 347912 5578
rect 348160 2990 348188 331214
rect 348436 15434 348464 335582
rect 348424 15428 348476 15434
rect 348424 15370 348476 15376
rect 349356 15298 349384 340054
rect 349448 336870 349476 340068
rect 349436 336864 349488 336870
rect 349436 336806 349488 336812
rect 349724 336802 349752 340068
rect 349712 336796 349764 336802
rect 349712 336738 349764 336744
rect 349816 22098 349844 459326
rect 349908 405686 349936 459410
rect 349896 405680 349948 405686
rect 349896 405622 349948 405628
rect 371882 310992 371938 311001
rect 371882 310927 371938 310936
rect 350446 310720 350502 310729
rect 350446 310655 350502 310664
rect 367006 310720 367062 310729
rect 367006 310655 367062 310664
rect 350460 310570 350488 310655
rect 350630 310584 350686 310593
rect 350460 310542 350630 310570
rect 350630 310519 350686 310528
rect 367020 310321 367048 310655
rect 371896 310593 371924 310927
rect 371882 310584 371938 310593
rect 371882 310519 371938 310528
rect 367006 310312 367062 310321
rect 367006 310247 367062 310256
rect 371882 264072 371938 264081
rect 371882 264007 371938 264016
rect 350446 263800 350502 263809
rect 350446 263735 350502 263744
rect 367006 263800 367062 263809
rect 367006 263735 367062 263744
rect 350460 263650 350488 263735
rect 350630 263664 350686 263673
rect 350460 263622 350630 263650
rect 350630 263599 350686 263608
rect 367020 263401 367048 263735
rect 371896 263673 371924 264007
rect 371882 263664 371938 263673
rect 371882 263599 371938 263608
rect 367006 263392 367062 263401
rect 367006 263327 367062 263336
rect 371882 217152 371938 217161
rect 371882 217087 371938 217096
rect 350446 216880 350502 216889
rect 350446 216815 350502 216824
rect 367006 216880 367062 216889
rect 367006 216815 367062 216824
rect 350460 216730 350488 216815
rect 350630 216744 350686 216753
rect 350460 216702 350630 216730
rect 350630 216679 350686 216688
rect 367020 216481 367048 216815
rect 371896 216753 371924 217087
rect 371882 216744 371938 216753
rect 371882 216679 371938 216688
rect 367006 216472 367062 216481
rect 367006 216407 367062 216416
rect 371882 170232 371938 170241
rect 371882 170167 371938 170176
rect 350446 169960 350502 169969
rect 350446 169895 350502 169904
rect 367006 169960 367062 169969
rect 367006 169895 367062 169904
rect 350460 169810 350488 169895
rect 350630 169824 350686 169833
rect 350460 169782 350630 169810
rect 350630 169759 350686 169768
rect 367020 169561 367048 169895
rect 371896 169833 371924 170167
rect 371882 169824 371938 169833
rect 371882 169759 371938 169768
rect 367006 169552 367062 169561
rect 367006 169487 367062 169496
rect 577516 124166 577544 462470
rect 580356 462460 580408 462466
rect 580356 462402 580408 462408
rect 580172 460284 580224 460290
rect 580172 460226 580224 460232
rect 579988 460012 580040 460018
rect 579988 459954 580040 459960
rect 579712 459876 579764 459882
rect 579712 459818 579764 459824
rect 579724 451654 579752 459818
rect 579896 459128 579948 459134
rect 579896 459070 579948 459076
rect 579802 457872 579858 457881
rect 579802 457807 579858 457816
rect 579712 451648 579764 451654
rect 579712 451590 579764 451596
rect 579816 439929 579844 457807
rect 579802 439920 579858 439929
rect 579802 439855 579858 439864
rect 579804 405680 579856 405686
rect 579804 405622 579856 405628
rect 579816 404841 579844 405622
rect 579802 404832 579858 404841
rect 579802 404767 579858 404776
rect 579908 357921 579936 459070
rect 579894 357912 579950 357921
rect 579894 357847 579950 357856
rect 580000 322697 580028 459954
rect 580080 458856 580132 458862
rect 580080 458798 580132 458804
rect 579986 322688 580042 322697
rect 579986 322623 580042 322632
rect 580092 299169 580120 458798
rect 580184 451761 580212 460226
rect 580264 459604 580316 459610
rect 580264 459546 580316 459552
rect 580170 451752 580226 451761
rect 580170 451687 580226 451696
rect 580172 451648 580224 451654
rect 580172 451590 580224 451596
rect 580078 299160 580134 299169
rect 580078 299095 580134 299104
rect 580184 275777 580212 451590
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 577504 124160 577556 124166
rect 577504 124102 577556 124108
rect 579620 124160 579672 124166
rect 579620 124102 579672 124108
rect 579632 123185 579660 124102
rect 579618 123176 579674 123185
rect 579618 123111 579674 123120
rect 375286 87408 375342 87417
rect 375286 87343 375342 87352
rect 350446 87136 350502 87145
rect 360290 87136 360346 87145
rect 350502 87094 350672 87122
rect 350446 87071 350502 87080
rect 350644 87009 350672 87094
rect 360290 87071 360346 87080
rect 350630 87000 350686 87009
rect 350630 86935 350686 86944
rect 360106 87000 360162 87009
rect 360304 86986 360332 87071
rect 375300 87009 375328 87343
rect 386326 87272 386382 87281
rect 386326 87207 386382 87216
rect 386340 87174 386368 87207
rect 379428 87168 379480 87174
rect 379426 87136 379428 87145
rect 386328 87168 386380 87174
rect 379480 87136 379482 87145
rect 386328 87110 386380 87116
rect 379426 87071 379482 87080
rect 360162 86958 360332 86986
rect 375286 87000 375342 87009
rect 360106 86935 360162 86944
rect 375286 86935 375342 86944
rect 580276 76265 580304 459546
rect 580368 111489 580396 462402
rect 580816 459740 580868 459746
rect 580816 459682 580868 459688
rect 580632 459672 580684 459678
rect 580632 459614 580684 459620
rect 580540 458312 580592 458318
rect 580540 458254 580592 458260
rect 580448 458244 580500 458250
rect 580448 458186 580500 458192
rect 580460 134881 580488 458186
rect 580552 158409 580580 458254
rect 580644 181937 580672 459614
rect 580724 458516 580776 458522
rect 580724 458458 580776 458464
rect 580736 205329 580764 458458
rect 580828 228857 580856 459682
rect 580908 458584 580960 458590
rect 580908 458526 580960 458532
rect 580920 252249 580948 458526
rect 580906 252240 580962 252249
rect 580906 252175 580962 252184
rect 580814 228848 580870 228857
rect 580814 228783 580870 228792
rect 580722 205320 580778 205329
rect 580722 205255 580778 205264
rect 580630 181928 580686 181937
rect 580630 181863 580686 181872
rect 580538 158400 580594 158409
rect 580538 158335 580594 158344
rect 580446 134872 580502 134881
rect 580446 134807 580502 134816
rect 580354 111480 580410 111489
rect 580354 111415 580410 111424
rect 580262 76256 580318 76265
rect 580262 76191 580318 76200
rect 353206 64016 353262 64025
rect 353206 63951 353262 63960
rect 371882 64016 371938 64025
rect 371882 63951 371938 63960
rect 353220 63753 353248 63951
rect 353206 63744 353262 63753
rect 353206 63679 353262 63688
rect 354586 63744 354642 63753
rect 354586 63679 354642 63688
rect 367006 63744 367062 63753
rect 367006 63679 367062 63688
rect 354600 63617 354628 63679
rect 354586 63608 354642 63617
rect 354586 63543 354642 63552
rect 364246 63472 364302 63481
rect 364246 63407 364302 63416
rect 364260 63345 364288 63407
rect 367020 63345 367048 63679
rect 371896 63617 371924 63951
rect 371882 63608 371938 63617
rect 371882 63543 371938 63552
rect 364246 63336 364302 63345
rect 364246 63271 364302 63280
rect 367006 63336 367062 63345
rect 367006 63271 367062 63280
rect 355966 40624 356022 40633
rect 355966 40559 356022 40568
rect 355980 40089 356008 40559
rect 371882 40488 371938 40497
rect 371882 40423 371938 40432
rect 367006 40216 367062 40225
rect 367006 40151 367062 40160
rect 355966 40080 356022 40089
rect 355966 40015 356022 40024
rect 367020 39817 367048 40151
rect 371896 40089 371924 40423
rect 371882 40080 371938 40089
rect 371882 40015 371938 40024
rect 367006 39808 367062 39817
rect 367006 39743 367062 39752
rect 355966 29472 356022 29481
rect 355966 29407 356022 29416
rect 375286 29472 375342 29481
rect 375286 29407 375342 29416
rect 355980 29073 356008 29407
rect 360290 29200 360346 29209
rect 360120 29158 360290 29186
rect 360120 29073 360148 29158
rect 360290 29135 360346 29144
rect 375300 29073 375328 29407
rect 386326 29336 386382 29345
rect 386326 29271 386382 29280
rect 386340 29238 386368 29271
rect 379428 29232 379480 29238
rect 379426 29200 379428 29209
rect 386328 29232 386380 29238
rect 379480 29200 379482 29209
rect 386328 29174 386380 29180
rect 379426 29135 379482 29144
rect 355966 29064 356022 29073
rect 355966 28999 356022 29008
rect 360106 29064 360162 29073
rect 360106 28999 360162 29008
rect 375286 29064 375342 29073
rect 375286 28999 375342 29008
rect 349804 22092 349856 22098
rect 349804 22034 349856 22040
rect 443000 18556 443052 18562
rect 443000 18498 443052 18504
rect 431960 17944 432012 17950
rect 431960 17886 432012 17892
rect 390560 17196 390612 17202
rect 390560 17138 390612 17144
rect 387800 17128 387852 17134
rect 387800 17070 387852 17076
rect 369766 16824 369822 16833
rect 379610 16824 379666 16833
rect 369766 16759 369822 16768
rect 379440 16782 379610 16810
rect 369780 16674 369808 16759
rect 379440 16697 379468 16782
rect 379610 16759 379666 16768
rect 369950 16688 370006 16697
rect 369780 16646 369950 16674
rect 369950 16623 370006 16632
rect 379426 16688 379482 16697
rect 379426 16623 379482 16632
rect 349344 15292 349396 15298
rect 349344 15234 349396 15240
rect 374000 13796 374052 13802
rect 374000 13738 374052 13744
rect 371240 13048 371292 13054
rect 371240 12990 371292 12996
rect 367100 12980 367152 12986
rect 367100 12922 367152 12928
rect 364340 12912 364392 12918
rect 364340 12854 364392 12860
rect 360200 12844 360252 12850
rect 360200 12786 360252 12792
rect 356060 12776 356112 12782
rect 356060 12718 356112 12724
rect 353300 12708 353352 12714
rect 353300 12650 353352 12656
rect 349160 12640 349212 12646
rect 349160 12582 349212 12588
rect 349068 8764 349120 8770
rect 349068 8706 349120 8712
rect 348148 2984 348200 2990
rect 348148 2926 348200 2932
rect 349080 480 349108 8706
rect 349172 610 349200 12582
rect 352564 8832 352616 8838
rect 352564 8774 352616 8780
rect 351368 5704 351420 5710
rect 351368 5646 351420 5652
rect 349160 604 349212 610
rect 349160 546 349212 552
rect 350264 604 350316 610
rect 350264 546 350316 552
rect 350276 480 350304 546
rect 351380 480 351408 5646
rect 352576 480 352604 8774
rect 353312 626 353340 12650
rect 354956 5772 355008 5778
rect 354956 5714 355008 5720
rect 353312 598 353800 626
rect 353772 480 353800 598
rect 354968 480 354996 5714
rect 356072 882 356100 12718
rect 359740 9648 359792 9654
rect 359740 9590 359792 9596
rect 356152 8900 356204 8906
rect 356152 8842 356204 8848
rect 356060 876 356112 882
rect 356060 818 356112 824
rect 356164 480 356192 8842
rect 358544 5840 358596 5846
rect 358544 5782 358596 5788
rect 357348 876 357400 882
rect 357348 818 357400 824
rect 357360 480 357388 818
rect 358556 480 358584 5782
rect 359752 480 359780 9590
rect 360212 3346 360240 12786
rect 363328 9580 363380 9586
rect 363328 9522 363380 9528
rect 362132 5908 362184 5914
rect 362132 5850 362184 5856
rect 360212 3318 360976 3346
rect 360948 480 360976 3318
rect 362144 480 362172 5850
rect 363340 480 363368 9522
rect 364352 3346 364380 12854
rect 366916 9512 366968 9518
rect 366916 9454 366968 9460
rect 365720 5976 365772 5982
rect 365720 5918 365772 5924
rect 364352 3318 364564 3346
rect 364536 480 364564 3318
rect 365732 480 365760 5918
rect 366928 480 366956 9454
rect 367112 3346 367140 12922
rect 370412 9444 370464 9450
rect 370412 9386 370464 9392
rect 369216 6044 369268 6050
rect 369216 5986 369268 5992
rect 367112 3318 368060 3346
rect 368032 480 368060 3318
rect 369228 480 369256 5986
rect 370424 480 370452 9386
rect 371252 3346 371280 12990
rect 372804 6112 372856 6118
rect 372804 6054 372856 6060
rect 371252 3318 371648 3346
rect 371620 480 371648 3318
rect 372816 480 372844 6054
rect 374012 3398 374040 13738
rect 378140 13728 378192 13734
rect 378140 13670 378192 13676
rect 374092 9376 374144 9382
rect 374092 9318 374144 9324
rect 374000 3392 374052 3398
rect 374000 3334 374052 3340
rect 374104 1442 374132 9318
rect 377588 9308 377640 9314
rect 377588 9250 377640 9256
rect 376392 6860 376444 6866
rect 376392 6802 376444 6808
rect 375196 3392 375248 3398
rect 375196 3334 375248 3340
rect 374012 1414 374132 1442
rect 374012 480 374040 1414
rect 375208 480 375236 3334
rect 376404 480 376432 6802
rect 377600 480 377628 9250
rect 378152 3346 378180 13670
rect 382280 13660 382332 13666
rect 382280 13602 382332 13608
rect 381176 9240 381228 9246
rect 381176 9182 381228 9188
rect 379980 6792 380032 6798
rect 379980 6734 380032 6740
rect 378152 3318 378824 3346
rect 378796 480 378824 3318
rect 379992 480 380020 6734
rect 381188 480 381216 9182
rect 382292 3482 382320 13602
rect 385040 13592 385092 13598
rect 385040 13534 385092 13540
rect 384670 9616 384726 9625
rect 384670 9551 384726 9560
rect 383568 6724 383620 6730
rect 383568 6666 383620 6672
rect 382292 3454 382412 3482
rect 382384 480 382412 3454
rect 383580 480 383608 6666
rect 384684 480 384712 9551
rect 385052 3346 385080 13534
rect 387064 6656 387116 6662
rect 387064 6598 387116 6604
rect 385052 3318 385908 3346
rect 385880 480 385908 3318
rect 387076 480 387104 6598
rect 387812 3346 387840 17070
rect 389086 16824 389142 16833
rect 389142 16782 389312 16810
rect 389086 16759 389142 16768
rect 389284 16697 389312 16782
rect 389270 16688 389326 16697
rect 389270 16623 389326 16632
rect 389180 13524 389232 13530
rect 389180 13466 389232 13472
rect 389192 3346 389220 13466
rect 390572 3398 390600 17138
rect 404266 16824 404322 16833
rect 404266 16759 404322 16768
rect 408406 16824 408462 16833
rect 408406 16759 408462 16768
rect 404280 16726 404308 16759
rect 394700 16720 394752 16726
rect 394698 16688 394700 16697
rect 404268 16720 404320 16726
rect 394752 16688 394754 16697
rect 404268 16662 404320 16668
rect 408420 16674 408448 16759
rect 408590 16688 408646 16697
rect 408420 16646 408590 16674
rect 394698 16623 394754 16632
rect 408590 16623 408646 16632
rect 414018 13696 414074 13705
rect 414018 13631 414074 13640
rect 391940 13456 391992 13462
rect 391940 13398 391992 13404
rect 390652 6588 390704 6594
rect 390652 6530 390704 6536
rect 390560 3392 390612 3398
rect 387812 3318 388300 3346
rect 389192 3318 389496 3346
rect 390560 3334 390612 3340
rect 388272 480 388300 3318
rect 389468 480 389496 3318
rect 390664 480 390692 6530
rect 391848 3392 391900 3398
rect 391848 3334 391900 3340
rect 391952 3346 391980 13398
rect 396080 13388 396132 13394
rect 396080 13330 396132 13336
rect 394700 9716 394752 9722
rect 394700 9658 394752 9664
rect 394240 6520 394292 6526
rect 394240 6462 394292 6468
rect 391860 480 391888 3334
rect 391952 3318 393084 3346
rect 393056 480 393084 3318
rect 394252 480 394280 6462
rect 394712 610 394740 9658
rect 396092 626 396120 13330
rect 400220 13320 400272 13326
rect 400220 13262 400272 13268
rect 398840 9784 398892 9790
rect 398840 9726 398892 9732
rect 397828 6452 397880 6458
rect 397828 6394 397880 6400
rect 394700 604 394752 610
rect 394700 546 394752 552
rect 395436 604 395488 610
rect 396092 598 396580 626
rect 396552 592 396580 598
rect 396552 564 396672 592
rect 395436 546 395488 552
rect 395448 480 395476 546
rect 396644 480 396672 564
rect 397840 480 397868 6394
rect 398852 626 398880 9726
rect 398852 598 398972 626
rect 398944 592 398972 598
rect 398944 564 399064 592
rect 399036 480 399064 564
rect 400232 480 400260 13262
rect 402980 13252 403032 13258
rect 402980 13194 403032 13200
rect 401600 9852 401652 9858
rect 401600 9794 401652 9800
rect 401324 6384 401376 6390
rect 401324 6326 401376 6332
rect 401336 480 401364 6326
rect 401612 610 401640 9794
rect 402992 610 403020 13194
rect 407120 13184 407172 13190
rect 407120 13126 407172 13132
rect 405740 9920 405792 9926
rect 405740 9862 405792 9868
rect 404912 6316 404964 6322
rect 404912 6258 404964 6264
rect 401600 604 401652 610
rect 401600 546 401652 552
rect 402520 604 402572 610
rect 402520 546 402572 552
rect 402980 604 403032 610
rect 402980 546 403032 552
rect 403716 604 403768 610
rect 403716 546 403768 552
rect 402532 480 402560 546
rect 403728 480 403756 546
rect 404924 480 404952 6258
rect 405752 610 405780 9862
rect 407132 626 407160 13126
rect 409880 13116 409932 13122
rect 409880 13058 409932 13064
rect 408500 9988 408552 9994
rect 408500 9930 408552 9936
rect 408512 3398 408540 9930
rect 408592 6248 408644 6254
rect 408592 6190 408644 6196
rect 408500 3392 408552 3398
rect 408500 3334 408552 3340
rect 408604 3210 408632 6190
rect 409696 3392 409748 3398
rect 409696 3334 409748 3340
rect 408512 3182 408632 3210
rect 405740 604 405792 610
rect 405740 546 405792 552
rect 406108 604 406160 610
rect 407132 598 407344 626
rect 406108 546 406160 552
rect 406120 480 406148 546
rect 407316 480 407344 598
rect 408512 480 408540 3182
rect 409708 480 409736 3334
rect 409892 610 409920 13058
rect 412640 10056 412692 10062
rect 412640 9998 412692 10004
rect 412088 6180 412140 6186
rect 412088 6122 412140 6128
rect 409880 604 409932 610
rect 409880 546 409932 552
rect 410892 604 410944 610
rect 410892 546 410944 552
rect 410904 480 410932 546
rect 412100 480 412128 6122
rect 412652 3346 412680 9998
rect 414032 3346 414060 13631
rect 416778 13560 416834 13569
rect 416778 13495 416834 13504
rect 415674 6760 415730 6769
rect 415674 6695 415730 6704
rect 412652 3318 413324 3346
rect 414032 3318 414520 3346
rect 413296 480 413324 3318
rect 414492 480 414520 3318
rect 415688 480 415716 6695
rect 416792 3398 416820 13495
rect 420918 13424 420974 13433
rect 420918 13359 420974 13368
rect 419540 10192 419592 10198
rect 419540 10134 419592 10140
rect 416872 10124 416924 10130
rect 416872 10066 416924 10072
rect 416780 3392 416832 3398
rect 416780 3334 416832 3340
rect 416884 480 416912 10066
rect 419170 6624 419226 6633
rect 419170 6559 419226 6568
rect 417976 3392 418028 3398
rect 417976 3334 418028 3340
rect 417988 480 418016 3334
rect 419184 480 419212 6559
rect 419552 3346 419580 10134
rect 420932 3346 420960 13359
rect 425058 13288 425114 13297
rect 425058 13223 425114 13232
rect 423680 10260 423732 10266
rect 423680 10202 423732 10208
rect 422758 6488 422814 6497
rect 422758 6423 422814 6432
rect 419552 3318 420408 3346
rect 420932 3318 421604 3346
rect 420380 480 420408 3318
rect 421576 480 421604 3318
rect 422772 480 422800 6423
rect 423692 610 423720 10202
rect 425072 626 425100 13223
rect 427818 13152 427874 13161
rect 427818 13087 427874 13096
rect 426440 11008 426492 11014
rect 426440 10950 426492 10956
rect 426346 6352 426402 6361
rect 426346 6287 426402 6296
rect 423680 604 423732 610
rect 423680 546 423732 552
rect 423956 604 424008 610
rect 425072 598 425192 626
rect 423956 546 424008 552
rect 423968 480 423996 546
rect 425164 480 425192 598
rect 426360 480 426388 6287
rect 426452 610 426480 10950
rect 427832 610 427860 13087
rect 430580 10940 430632 10946
rect 430580 10882 430632 10888
rect 429934 6216 429990 6225
rect 429934 6151 429990 6160
rect 426440 604 426492 610
rect 426440 546 426492 552
rect 427544 604 427596 610
rect 427544 546 427596 552
rect 427820 604 427872 610
rect 427820 546 427872 552
rect 428740 604 428792 610
rect 428740 546 428792 552
rect 427556 480 427584 546
rect 428752 480 428780 546
rect 429948 480 429976 6151
rect 430592 610 430620 10882
rect 431972 626 432000 17886
rect 433340 17876 433392 17882
rect 433340 17818 433392 17824
rect 433352 3482 433380 17818
rect 434720 17808 434772 17814
rect 434720 17750 434772 17756
rect 433432 10872 433484 10878
rect 433432 10814 433484 10820
rect 433444 3670 433472 10814
rect 433432 3664 433484 3670
rect 433432 3606 433484 3612
rect 434628 3664 434680 3670
rect 434628 3606 434680 3612
rect 433352 3454 433564 3482
rect 430580 604 430632 610
rect 430580 546 430632 552
rect 431132 604 431184 610
rect 431972 598 432368 626
rect 431132 546 431184 552
rect 431144 480 431172 546
rect 432340 480 432368 598
rect 433536 480 433564 3454
rect 434640 480 434668 3606
rect 434732 610 434760 17750
rect 436100 17740 436152 17746
rect 436100 17682 436152 17688
rect 436112 610 436140 17682
rect 438860 17672 438912 17678
rect 438860 17614 438912 17620
rect 437386 16688 437442 16697
rect 437386 16623 437388 16632
rect 437440 16623 437442 16632
rect 437388 16594 437440 16600
rect 437480 10804 437532 10810
rect 437480 10746 437532 10752
rect 437492 610 437520 10746
rect 438872 610 438900 17614
rect 440240 17604 440292 17610
rect 440240 17546 440292 17552
rect 440252 626 440280 17546
rect 442906 16688 442962 16697
rect 442906 16623 442908 16632
rect 442960 16623 442962 16632
rect 442908 16594 442960 16600
rect 441620 10736 441672 10742
rect 441620 10678 441672 10684
rect 441632 3482 441660 10678
rect 441632 3454 441844 3482
rect 434720 604 434772 610
rect 434720 546 434772 552
rect 435824 604 435876 610
rect 435824 546 435876 552
rect 436100 604 436152 610
rect 436100 546 436152 552
rect 437020 604 437072 610
rect 437020 546 437072 552
rect 437480 604 437532 610
rect 437480 546 437532 552
rect 438216 604 438268 610
rect 438216 546 438268 552
rect 438860 604 438912 610
rect 438860 546 438912 552
rect 439412 604 439464 610
rect 440252 598 440648 626
rect 439412 546 439464 552
rect 435836 480 435864 546
rect 437032 480 437060 546
rect 438228 480 438256 546
rect 439424 480 439452 546
rect 440620 480 440648 598
rect 441816 480 441844 3454
rect 443012 480 443040 18498
rect 492678 17776 492734 17785
rect 492678 17711 492734 17720
rect 483020 17536 483072 17542
rect 483020 17478 483072 17484
rect 447046 16824 447102 16833
rect 447230 16824 447286 16833
rect 447102 16782 447230 16810
rect 447046 16759 447102 16768
rect 447230 16759 447286 16768
rect 466366 16824 466422 16833
rect 476210 16824 476266 16833
rect 466366 16759 466422 16768
rect 476040 16782 476210 16810
rect 466380 16674 466408 16759
rect 476040 16697 476068 16782
rect 476210 16759 476266 16768
rect 466550 16688 466606 16697
rect 466380 16646 466550 16674
rect 466550 16623 466606 16632
rect 476026 16688 476082 16697
rect 476026 16623 476082 16632
rect 477500 15156 477552 15162
rect 477500 15098 477552 15104
rect 474740 14408 474792 14414
rect 474740 14350 474792 14356
rect 470600 14340 470652 14346
rect 470600 14282 470652 14288
rect 467840 14272 467892 14278
rect 467840 14214 467892 14220
rect 463700 14204 463752 14210
rect 463700 14146 463752 14152
rect 459560 14136 459612 14142
rect 459560 14078 459612 14084
rect 456800 14068 456852 14074
rect 456800 14010 456852 14016
rect 452660 14000 452712 14006
rect 452660 13942 452712 13948
rect 449900 13932 449952 13938
rect 449900 13874 449952 13880
rect 445760 13864 445812 13870
rect 445760 13806 445812 13812
rect 444380 10668 444432 10674
rect 444380 10610 444432 10616
rect 444196 7064 444248 7070
rect 444196 7006 444248 7012
rect 444208 480 444236 7006
rect 444392 3482 444420 10610
rect 445772 3482 445800 13806
rect 448520 10600 448572 10606
rect 448520 10542 448572 10548
rect 447784 7132 447836 7138
rect 447784 7074 447836 7080
rect 444392 3454 445432 3482
rect 445772 3454 446628 3482
rect 445404 480 445432 3454
rect 446600 480 446628 3454
rect 447796 480 447824 7074
rect 448532 3482 448560 10542
rect 449912 3482 449940 13874
rect 451280 10532 451332 10538
rect 451280 10474 451332 10480
rect 448532 3454 449020 3482
rect 449912 3454 450216 3482
rect 448992 480 449020 3454
rect 450188 480 450216 3454
rect 451292 3398 451320 10474
rect 451372 7200 451424 7206
rect 451372 7142 451424 7148
rect 451280 3392 451332 3398
rect 451280 3334 451332 3340
rect 451384 1442 451412 7142
rect 452476 3392 452528 3398
rect 452476 3334 452528 3340
rect 451292 1414 451412 1442
rect 451292 480 451320 1414
rect 452488 480 452516 3334
rect 452672 610 452700 13942
rect 455420 10464 455472 10470
rect 455420 10406 455472 10412
rect 454868 7268 454920 7274
rect 454868 7210 454920 7216
rect 452660 604 452712 610
rect 452660 546 452712 552
rect 453672 604 453724 610
rect 453672 546 453724 552
rect 453684 480 453712 546
rect 454880 480 454908 7210
rect 455432 610 455460 10406
rect 456812 610 456840 14010
rect 458456 7336 458508 7342
rect 458456 7278 458508 7284
rect 455420 604 455472 610
rect 455420 546 455472 552
rect 456064 604 456116 610
rect 456064 546 456116 552
rect 456800 604 456852 610
rect 456800 546 456852 552
rect 457260 604 457312 610
rect 457260 546 457312 552
rect 456076 480 456104 546
rect 457272 480 457300 546
rect 458468 480 458496 7278
rect 459572 3398 459600 14078
rect 459652 10396 459704 10402
rect 459652 10338 459704 10344
rect 459560 3392 459612 3398
rect 459560 3334 459612 3340
rect 459664 480 459692 10338
rect 462320 10328 462372 10334
rect 462320 10270 462372 10276
rect 462044 7404 462096 7410
rect 462044 7346 462096 7352
rect 460848 3392 460900 3398
rect 460848 3334 460900 3340
rect 460860 480 460888 3334
rect 462056 480 462084 7346
rect 462332 610 462360 10270
rect 463712 610 463740 14146
rect 466458 10840 466514 10849
rect 466458 10775 466514 10784
rect 465632 7472 465684 7478
rect 465632 7414 465684 7420
rect 462320 604 462372 610
rect 462320 546 462372 552
rect 463240 604 463292 610
rect 463240 546 463292 552
rect 463700 604 463752 610
rect 463700 546 463752 552
rect 464436 604 464488 610
rect 464436 546 464488 552
rect 463252 480 463280 546
rect 464448 480 464476 546
rect 465644 480 465672 7414
rect 466472 610 466500 10775
rect 467852 626 467880 14214
rect 469218 10704 469274 10713
rect 469218 10639 469274 10648
rect 469128 7540 469180 7546
rect 469128 7482 469180 7488
rect 466460 604 466512 610
rect 466460 546 466512 552
rect 466828 604 466880 610
rect 467852 598 467972 626
rect 466828 546 466880 552
rect 466840 480 466868 546
rect 467944 480 467972 598
rect 469140 480 469168 7482
rect 469232 610 469260 10639
rect 470612 610 470640 14282
rect 473358 10568 473414 10577
rect 473358 10503 473414 10512
rect 472716 8288 472768 8294
rect 472716 8230 472768 8236
rect 469220 604 469272 610
rect 469220 546 469272 552
rect 470324 604 470376 610
rect 470324 546 470376 552
rect 470600 604 470652 610
rect 470600 546 470652 552
rect 471520 604 471572 610
rect 471520 546 471572 552
rect 470336 480 470364 546
rect 471532 480 471560 546
rect 472728 480 472756 8230
rect 473372 626 473400 10503
rect 474752 626 474780 14350
rect 476304 8220 476356 8226
rect 476304 8162 476356 8168
rect 473372 598 473860 626
rect 474752 598 475056 626
rect 473832 592 473860 598
rect 475028 592 475056 598
rect 473832 564 473952 592
rect 475028 564 475148 592
rect 473924 480 473952 564
rect 475120 480 475148 564
rect 476316 480 476344 8162
rect 477512 3670 477540 15098
rect 481640 15088 481692 15094
rect 481640 15030 481692 15036
rect 477590 10432 477646 10441
rect 477590 10367 477646 10376
rect 477500 3664 477552 3670
rect 477500 3606 477552 3612
rect 477604 3482 477632 10367
rect 480258 10296 480314 10305
rect 480258 10231 480314 10240
rect 479892 8152 479944 8158
rect 479892 8094 479944 8100
rect 478696 3664 478748 3670
rect 478696 3606 478748 3612
rect 477512 3454 477632 3482
rect 477512 480 477540 3454
rect 478708 480 478736 3606
rect 479904 480 479932 8094
rect 480272 3482 480300 10231
rect 481652 3482 481680 15030
rect 483032 3482 483060 17478
rect 485780 17468 485832 17474
rect 485780 17410 485832 17416
rect 484584 8084 484636 8090
rect 484584 8026 484636 8032
rect 480272 3454 481128 3482
rect 481652 3454 482324 3482
rect 483032 3454 483520 3482
rect 481100 480 481128 3454
rect 482296 480 482324 3454
rect 483492 480 483520 3454
rect 484596 480 484624 8026
rect 485792 3670 485820 17410
rect 485872 17400 485924 17406
rect 485872 17342 485924 17348
rect 485780 3664 485832 3670
rect 485780 3606 485832 3612
rect 485884 3482 485912 17342
rect 488540 17332 488592 17338
rect 488540 17274 488592 17280
rect 488172 8016 488224 8022
rect 488172 7958 488224 7964
rect 486976 3664 487028 3670
rect 486976 3606 487028 3612
rect 485792 3454 485912 3482
rect 485792 480 485820 3454
rect 486988 480 487016 3606
rect 488184 480 488212 7958
rect 488552 3482 488580 17274
rect 489920 17264 489972 17270
rect 489920 17206 489972 17212
rect 488552 3454 489408 3482
rect 489380 480 489408 3454
rect 489932 610 489960 17206
rect 491206 16824 491262 16833
rect 491206 16759 491262 16768
rect 491220 16561 491248 16759
rect 491206 16552 491262 16561
rect 491206 16487 491262 16496
rect 491760 7948 491812 7954
rect 491760 7890 491812 7896
rect 489920 604 489972 610
rect 489920 546 489972 552
rect 490564 604 490616 610
rect 490564 546 490616 552
rect 490576 480 490604 546
rect 491772 480 491800 7890
rect 492692 626 492720 17711
rect 534078 17640 534134 17649
rect 534078 17575 534134 17584
rect 495346 17096 495402 17105
rect 495530 17096 495586 17105
rect 495402 17054 495530 17082
rect 495346 17031 495402 17040
rect 495530 17031 495586 17040
rect 505006 16960 505062 16969
rect 505006 16895 505008 16904
rect 505060 16895 505062 16904
rect 511908 16924 511960 16930
rect 505008 16866 505060 16872
rect 511908 16866 511960 16872
rect 511920 16833 511948 16866
rect 511906 16824 511962 16833
rect 511906 16759 511962 16768
rect 520280 12436 520332 12442
rect 520280 12378 520332 12384
rect 517520 11688 517572 11694
rect 517520 11630 517572 11636
rect 513380 11620 513432 11626
rect 513380 11562 513432 11568
rect 510620 11552 510672 11558
rect 510620 11494 510672 11500
rect 506480 11484 506532 11490
rect 506480 11426 506532 11432
rect 502340 11416 502392 11422
rect 502340 11358 502392 11364
rect 499580 11348 499632 11354
rect 499580 11290 499632 11296
rect 495440 11280 495492 11286
rect 495440 11222 495492 11228
rect 495348 7880 495400 7886
rect 495348 7822 495400 7828
rect 494152 4276 494204 4282
rect 494152 4218 494204 4224
rect 492692 598 492904 626
rect 492876 592 492904 598
rect 492876 564 492996 592
rect 492968 480 492996 564
rect 494164 480 494192 4218
rect 495360 480 495388 7822
rect 495452 610 495480 11222
rect 498936 7812 498988 7818
rect 498936 7754 498988 7760
rect 497740 4344 497792 4350
rect 497740 4286 497792 4292
rect 495440 604 495492 610
rect 495440 546 495492 552
rect 496544 604 496596 610
rect 496544 546 496596 552
rect 496556 480 496584 546
rect 497752 480 497780 4286
rect 498948 480 498976 7754
rect 499592 610 499620 11290
rect 501236 4412 501288 4418
rect 501236 4354 501288 4360
rect 499580 604 499632 610
rect 499580 546 499632 552
rect 500132 604 500184 610
rect 500132 546 500184 552
rect 500144 480 500172 546
rect 501248 480 501276 4354
rect 502352 3398 502380 11358
rect 502432 7744 502484 7750
rect 502432 7686 502484 7692
rect 502340 3392 502392 3398
rect 502340 3334 502392 3340
rect 502444 480 502472 7686
rect 506020 7676 506072 7682
rect 506020 7618 506072 7624
rect 504824 4480 504876 4486
rect 504824 4422 504876 4428
rect 503628 3392 503680 3398
rect 503628 3334 503680 3340
rect 503640 480 503668 3334
rect 504836 480 504864 4422
rect 506032 480 506060 7618
rect 506492 610 506520 11426
rect 509606 8256 509662 8265
rect 509606 8191 509662 8200
rect 508412 4548 508464 4554
rect 508412 4490 508464 4496
rect 506480 604 506532 610
rect 506480 546 506532 552
rect 507216 604 507268 610
rect 507216 546 507268 552
rect 507228 480 507256 546
rect 508424 480 508452 4490
rect 509620 480 509648 8191
rect 510632 610 510660 11494
rect 513194 8120 513250 8129
rect 513194 8055 513250 8064
rect 512000 4616 512052 4622
rect 512000 4558 512052 4564
rect 510620 604 510672 610
rect 510620 546 510672 552
rect 510804 604 510856 610
rect 510804 546 510856 552
rect 510816 480 510844 546
rect 512012 480 512040 4558
rect 513208 480 513236 8055
rect 513392 610 513420 11562
rect 516782 7984 516838 7993
rect 516782 7919 516838 7928
rect 515588 4684 515640 4690
rect 515588 4626 515640 4632
rect 513380 604 513432 610
rect 513380 546 513432 552
rect 514392 604 514444 610
rect 514392 546 514444 552
rect 514404 480 514432 546
rect 515600 480 515628 4626
rect 516796 480 516824 7919
rect 517532 626 517560 11630
rect 519084 4752 519136 4758
rect 519084 4694 519136 4700
rect 517532 598 517928 626
rect 517900 480 517928 598
rect 519096 480 519124 4694
rect 520292 3398 520320 12378
rect 524420 12368 524472 12374
rect 524420 12310 524472 12316
rect 523866 7848 523922 7857
rect 523866 7783 523922 7792
rect 520372 7608 520424 7614
rect 520372 7550 520424 7556
rect 520280 3392 520332 3398
rect 520280 3334 520332 3340
rect 520384 1442 520412 7550
rect 522672 5500 522724 5506
rect 522672 5442 522724 5448
rect 521476 3392 521528 3398
rect 521476 3334 521528 3340
rect 520292 1414 520412 1442
rect 520292 480 520320 1414
rect 521488 480 521516 3334
rect 522684 480 522712 5442
rect 523880 480 523908 7783
rect 524432 610 524460 12310
rect 528560 12300 528612 12306
rect 528560 12242 528612 12248
rect 527454 7712 527510 7721
rect 527454 7647 527510 7656
rect 526260 5432 526312 5438
rect 526260 5374 526312 5380
rect 524420 604 524472 610
rect 524420 546 524472 552
rect 525064 604 525116 610
rect 525064 546 525116 552
rect 525076 480 525104 546
rect 526272 480 526300 5374
rect 527468 480 527496 7647
rect 528572 3482 528600 12242
rect 531320 12232 531372 12238
rect 531320 12174 531372 12180
rect 531042 7576 531098 7585
rect 531042 7511 531098 7520
rect 529848 5364 529900 5370
rect 529848 5306 529900 5312
rect 528572 3454 528692 3482
rect 528664 480 528692 3454
rect 529860 480 529888 5306
rect 531056 480 531084 7511
rect 531332 3482 531360 12174
rect 533436 5296 533488 5302
rect 533436 5238 533488 5244
rect 531332 3454 532280 3482
rect 532252 480 532280 3454
rect 533448 480 533476 5238
rect 534092 3482 534120 17575
rect 536838 17504 536894 17513
rect 536838 17439 536894 17448
rect 535460 12164 535512 12170
rect 535460 12106 535512 12112
rect 535472 3482 535500 12106
rect 534092 3454 534580 3482
rect 535472 3454 535776 3482
rect 534552 480 534580 3454
rect 535748 480 535776 3454
rect 536852 3398 536880 17439
rect 540978 17368 541034 17377
rect 540978 17303 541034 17312
rect 538220 12096 538272 12102
rect 538220 12038 538272 12044
rect 536932 5228 536984 5234
rect 536932 5170 536984 5176
rect 536840 3392 536892 3398
rect 536840 3334 536892 3340
rect 536944 480 536972 5170
rect 538128 3392 538180 3398
rect 538128 3334 538180 3340
rect 538140 480 538168 3334
rect 538232 610 538260 12038
rect 540520 5160 540572 5166
rect 540520 5102 540572 5108
rect 538220 604 538272 610
rect 538220 546 538272 552
rect 539324 604 539376 610
rect 539324 546 539376 552
rect 539336 480 539364 546
rect 540532 480 540560 5102
rect 540992 610 541020 17303
rect 560298 12336 560354 12345
rect 560298 12271 560354 12280
rect 542360 12028 542412 12034
rect 542360 11970 542412 11976
rect 542372 610 542400 11970
rect 546500 11960 546552 11966
rect 546500 11902 546552 11908
rect 545304 9172 545356 9178
rect 545304 9114 545356 9120
rect 544108 5092 544160 5098
rect 544108 5034 544160 5040
rect 540980 604 541032 610
rect 540980 546 541032 552
rect 541716 604 541768 610
rect 541716 546 541768 552
rect 542360 604 542412 610
rect 542360 546 542412 552
rect 542912 604 542964 610
rect 542912 546 542964 552
rect 541728 480 541756 546
rect 542924 480 542952 546
rect 544120 480 544148 5034
rect 545316 480 545344 9114
rect 546512 480 546540 11902
rect 549260 11892 549312 11898
rect 549260 11834 549312 11840
rect 548890 9480 548946 9489
rect 548890 9415 548946 9424
rect 547696 5024 547748 5030
rect 547696 4966 547748 4972
rect 547708 480 547736 4966
rect 548904 480 548932 9415
rect 549272 610 549300 11834
rect 553400 11824 553452 11830
rect 553400 11766 553452 11772
rect 552388 9104 552440 9110
rect 552388 9046 552440 9052
rect 551192 4956 551244 4962
rect 551192 4898 551244 4904
rect 549260 604 549312 610
rect 549260 546 549312 552
rect 550088 604 550140 610
rect 550088 546 550140 552
rect 550100 480 550128 546
rect 551204 480 551232 4898
rect 552400 480 552428 9046
rect 553412 626 553440 11766
rect 556160 11756 556212 11762
rect 556160 11698 556212 11704
rect 555974 9344 556030 9353
rect 555974 9279 556030 9288
rect 554780 4888 554832 4894
rect 554780 4830 554832 4836
rect 553412 598 553624 626
rect 553596 480 553624 598
rect 554792 480 554820 4830
rect 555988 480 556016 9279
rect 556172 610 556200 11698
rect 559562 9208 559618 9217
rect 559562 9143 559618 9152
rect 558368 4820 558420 4826
rect 558368 4762 558420 4768
rect 556160 604 556212 610
rect 556160 546 556212 552
rect 557172 604 557224 610
rect 557172 546 557224 552
rect 557184 480 557212 546
rect 558380 480 558408 4762
rect 559576 480 559604 9143
rect 560312 3482 560340 12271
rect 563058 12200 563114 12209
rect 563058 12135 563114 12144
rect 561954 5536 562010 5545
rect 561954 5471 562010 5480
rect 560312 3454 560800 3482
rect 560772 480 560800 3454
rect 561968 480 561996 5471
rect 563072 2514 563100 12135
rect 567198 12064 567254 12073
rect 567198 11999 567254 12008
rect 563150 9072 563206 9081
rect 563150 9007 563206 9016
rect 563060 2508 563112 2514
rect 563060 2450 563112 2456
rect 563164 480 563192 9007
rect 565542 5400 565598 5409
rect 565542 5335 565598 5344
rect 564348 2508 564400 2514
rect 564348 2450 564400 2456
rect 564360 480 564388 2450
rect 565556 480 565584 5335
rect 566740 3596 566792 3602
rect 566740 3538 566792 3544
rect 566752 480 566780 3538
rect 567212 3482 567240 11999
rect 574098 11928 574154 11937
rect 574098 11863 574154 11872
rect 570234 8936 570290 8945
rect 570234 8871 570290 8880
rect 569038 5264 569094 5273
rect 569038 5199 569094 5208
rect 567212 3454 567884 3482
rect 567856 480 567884 3454
rect 569052 480 569080 5199
rect 570248 480 570276 8871
rect 572626 5128 572682 5137
rect 572626 5063 572682 5072
rect 571432 3528 571484 3534
rect 571432 3470 571484 3476
rect 571444 480 571472 3470
rect 572640 480 572668 5063
rect 574112 3482 574140 11863
rect 578238 11792 578294 11801
rect 578238 11727 578294 11736
rect 577412 9036 577464 9042
rect 577412 8978 577464 8984
rect 576214 4992 576270 5001
rect 576214 4927 576270 4936
rect 573824 3460 573876 3466
rect 574112 3454 575060 3482
rect 573824 3402 573876 3408
rect 573836 480 573864 3402
rect 575032 480 575060 3454
rect 576228 480 576256 4927
rect 577424 480 577452 8978
rect 578252 626 578280 11727
rect 580998 11656 581054 11665
rect 580998 11591 581054 11600
rect 579802 4856 579858 4865
rect 579802 4791 579858 4800
rect 578252 598 578648 626
rect 578620 480 578648 598
rect 579816 480 579844 4791
rect 581012 3534 581040 11591
rect 581092 8968 581144 8974
rect 581092 8910 581144 8916
rect 581000 3528 581052 3534
rect 581000 3470 581052 3476
rect 581104 1442 581132 8910
rect 582196 3528 582248 3534
rect 582196 3470 582248 3476
rect 581012 1414 581132 1442
rect 581012 480 581040 1414
rect 582208 480 582236 3470
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3514 682216 3570 682272
rect 3422 667956 3478 667992
rect 3422 667936 3424 667956
rect 3424 667936 3476 667956
rect 3476 667936 3478 667956
rect 3054 653520 3110 653576
rect 3422 624824 3478 624880
rect 3422 610408 3478 610464
rect 3238 595992 3294 596048
rect 3422 567296 3478 567352
rect 3146 553016 3202 553072
rect 3422 538600 3478 538656
rect 3422 509904 3478 509960
rect 3422 495508 3478 495544
rect 3422 495488 3424 495508
rect 3424 495488 3476 495508
rect 3476 495488 3478 495508
rect 3146 481072 3202 481128
rect 218978 540912 219034 540968
rect 219162 540912 219218 540968
rect 218978 531256 219034 531312
rect 219162 531256 219218 531312
rect 218794 521600 218850 521656
rect 218978 521600 219034 521656
rect 154302 463664 154358 463720
rect 154486 463664 154542 463720
rect 252466 462984 252522 463040
rect 2778 437996 2780 438016
rect 2780 437996 2832 438016
rect 2832 437996 2834 438016
rect 2778 437960 2834 437996
rect 2962 423680 3018 423736
rect 3054 394984 3110 395040
rect 3146 380568 3202 380624
rect 3330 457680 3386 457736
rect 3238 366152 3294 366208
rect 3330 337456 3386 337512
rect 2778 323040 2834 323096
rect 2778 280100 2780 280120
rect 2780 280100 2832 280120
rect 2832 280100 2834 280120
rect 2778 280064 2834 280100
rect 2778 265648 2834 265704
rect 2778 236952 2834 237008
rect 2778 222536 2834 222592
rect 2778 193840 2834 193896
rect 2778 179424 2834 179480
rect 2778 150728 2834 150784
rect 2778 136348 2780 136368
rect 2780 136348 2832 136368
rect 2832 136348 2834 136368
rect 2778 136312 2834 136348
rect 3330 107616 3386 107672
rect 3330 50904 3386 50960
rect 3330 50088 3386 50144
rect 2870 21392 2926 21448
rect 2686 11736 2742 11792
rect 1306 11600 1362 11656
rect 4066 308760 4122 308816
rect 3974 294344 4030 294400
rect 3882 251232 3938 251288
rect 3790 208120 3846 208176
rect 3698 165008 3754 165064
rect 22006 337592 22062 337648
rect 12346 337456 12402 337512
rect 10966 337320 11022 337376
rect 3606 122032 3662 122088
rect 3514 93200 3570 93256
rect 3514 80008 3570 80064
rect 3514 78920 3570 78976
rect 4066 15816 4122 15872
rect 3974 12960 4030 13016
rect 3422 7112 3478 7168
rect 9586 15952 9642 16008
rect 8206 14456 8262 14512
rect 21914 16360 21970 16416
rect 17866 16224 17922 16280
rect 13726 16088 13782 16144
rect 13634 14592 13690 14648
rect 6458 3304 6514 3360
rect 16026 3576 16082 3632
rect 14830 3440 14886 3496
rect 18326 3712 18382 3768
rect 251638 459992 251694 460048
rect 248326 459856 248382 459912
rect 255594 462712 255650 462768
rect 253478 462440 253534 462496
rect 256606 462576 256662 462632
rect 245382 459720 245438 459776
rect 580170 697992 580226 698048
rect 494886 686024 494942 686080
rect 494242 685888 494298 685944
rect 580170 686296 580226 686352
rect 580170 674600 580226 674656
rect 580170 651072 580226 651128
rect 580170 639376 580226 639432
rect 580170 627680 580226 627736
rect 580170 604152 580226 604208
rect 580170 592456 580226 592512
rect 493874 579672 493930 579728
rect 494058 579672 494114 579728
rect 580170 580760 580226 580816
rect 494150 560224 494206 560280
rect 494334 560224 494390 560280
rect 580170 557232 580226 557288
rect 580170 545536 580226 545592
rect 494150 540912 494206 540968
rect 494334 540912 494390 540968
rect 580170 533840 580226 533896
rect 494150 521600 494206 521656
rect 494334 521600 494390 521656
rect 542542 521600 542598 521656
rect 542726 521600 542782 521656
rect 559102 521600 559158 521656
rect 559286 521600 559342 521656
rect 580170 510312 580226 510368
rect 493966 502288 494022 502344
rect 494242 502324 494244 502344
rect 494244 502324 494296 502344
rect 494296 502324 494298 502344
rect 494242 502288 494298 502324
rect 542358 502288 542414 502344
rect 542634 502324 542636 502344
rect 542636 502324 542688 502344
rect 542688 502324 542690 502344
rect 542634 502288 542690 502324
rect 558918 502288 558974 502344
rect 559194 502324 559196 502344
rect 559196 502324 559248 502344
rect 559248 502324 559250 502344
rect 559194 502288 559250 502324
rect 580170 498616 580226 498672
rect 493966 492632 494022 492688
rect 494150 492632 494206 492688
rect 542358 492632 542414 492688
rect 542542 492652 542598 492688
rect 542542 492632 542544 492652
rect 542544 492632 542596 492652
rect 542596 492632 542598 492652
rect 558918 492632 558974 492688
rect 559102 492652 559158 492688
rect 559102 492632 559104 492652
rect 559104 492632 559156 492652
rect 559156 492632 559158 492652
rect 580170 486784 580226 486840
rect 580078 463392 580134 463448
rect 318706 462848 318762 462904
rect 231674 459584 231730 459640
rect 232686 459584 232742 459640
rect 233790 459584 233846 459640
rect 242254 459584 242310 459640
rect 343730 459584 343786 459640
rect 345294 459584 345350 459640
rect 37186 337728 37242 337784
rect 27526 16496 27582 16552
rect 24306 3984 24362 4040
rect 23110 3848 23166 3904
rect 48226 14728 48282 14784
rect 52366 14864 52422 14920
rect 56414 15000 56470 15056
rect 59266 15136 59322 15192
rect 71686 17176 71742 17232
rect 107474 278704 107530 278760
rect 107658 278704 107714 278760
rect 107474 259392 107530 259448
rect 107658 259392 107714 259448
rect 107474 241712 107530 241768
rect 107474 241576 107530 241632
rect 107474 240080 107530 240136
rect 107658 240080 107714 240136
rect 100666 231784 100722 231840
rect 100850 231784 100906 231840
rect 107474 220768 107530 220824
rect 107658 220768 107714 220824
rect 100666 212472 100722 212528
rect 100850 212472 100906 212528
rect 107474 211112 107530 211168
rect 107658 211112 107714 211168
rect 100666 193160 100722 193216
rect 100850 193160 100906 193216
rect 107474 191800 107530 191856
rect 107658 191800 107714 191856
rect 100666 173848 100722 173904
rect 100850 173848 100906 173904
rect 107474 172488 107530 172544
rect 107658 172488 107714 172544
rect 100666 164192 100722 164248
rect 100850 164192 100906 164248
rect 100666 144880 100722 144936
rect 100850 144880 100906 144936
rect 100666 125568 100722 125624
rect 100850 125568 100906 125624
rect 100482 9696 100538 9752
rect 100666 9696 100722 9752
rect 150438 8200 150494 8256
rect 146850 8064 146906 8120
rect 143262 7928 143318 7984
rect 139674 7792 139730 7848
rect 136086 7656 136142 7712
rect 132590 7520 132646 7576
rect 131394 6160 131450 6216
rect 130198 4800 130254 4856
rect 134890 6296 134946 6352
rect 138478 6432 138534 6488
rect 137282 4936 137338 4992
rect 142066 6568 142122 6624
rect 145654 6704 145710 6760
rect 149242 6840 149298 6896
rect 176566 5072 176622 5128
rect 183742 5208 183798 5264
rect 190826 5344 190882 5400
rect 234342 459312 234398 459368
rect 258814 459312 258870 459368
rect 324870 459312 324926 459368
rect 345754 459312 345810 459368
rect 347226 459312 347282 459368
rect 229098 16768 229154 16824
rect 205086 5480 205142 5536
rect 224774 3168 224830 3224
rect 224958 3168 225014 3224
rect 231214 338000 231270 338056
rect 230846 7520 230902 7576
rect 230754 6160 230810 6216
rect 231582 338000 231638 338056
rect 231766 258032 231822 258088
rect 231214 241440 231270 241496
rect 231398 241440 231454 241496
rect 231214 222128 231270 222184
rect 231398 222128 231454 222184
rect 231214 202816 231270 202872
rect 231398 202816 231454 202872
rect 231214 183504 231270 183560
rect 231398 183504 231454 183560
rect 231214 144880 231270 144936
rect 231398 144880 231454 144936
rect 231214 125568 231270 125624
rect 231398 125568 231454 125624
rect 231214 6296 231270 6352
rect 231950 278704 232006 278760
rect 232134 278704 232190 278760
rect 231950 258032 232006 258088
rect 232042 220768 232098 220824
rect 232042 211112 232098 211168
rect 232042 202816 232098 202872
rect 232134 202680 232190 202736
rect 232134 182144 232190 182200
rect 231950 172488 232006 172544
rect 232134 172488 232190 172544
rect 232318 240080 232374 240136
rect 232318 220768 232374 220824
rect 232318 182164 232374 182200
rect 232318 182144 232320 182164
rect 232320 182144 232372 182164
rect 232372 182144 232374 182164
rect 232594 240080 232650 240136
rect 232778 220768 232834 220824
rect 232502 139576 232558 139632
rect 232502 139440 232558 139496
rect 232318 7792 232374 7848
rect 232226 7656 232282 7712
rect 232042 6432 232098 6488
rect 232594 136584 232650 136640
rect 232870 136584 232926 136640
rect 232686 107616 232742 107672
rect 232870 107616 232926 107672
rect 232594 6568 232650 6624
rect 231858 4936 231914 4992
rect 233514 8064 233570 8120
rect 233422 7928 233478 7984
rect 233698 6704 233754 6760
rect 234894 8200 234950 8256
rect 234802 6840 234858 6896
rect 237838 240080 237894 240136
rect 238022 240080 238078 240136
rect 238666 90480 238722 90536
rect 238666 87080 238722 87136
rect 230570 4800 230626 4856
rect 240506 240080 240562 240136
rect 240506 220768 240562 220824
rect 240506 211112 240562 211168
rect 240690 240080 240746 240136
rect 240690 220768 240746 220824
rect 240690 211132 240746 211168
rect 240690 211112 240692 211132
rect 240692 211112 240744 211132
rect 240744 211112 240746 211132
rect 240690 201456 240746 201512
rect 240874 201456 240930 201512
rect 240690 182144 240746 182200
rect 240874 182144 240930 182200
rect 240690 162832 240746 162888
rect 240874 162832 240930 162888
rect 240690 143540 240746 143576
rect 240690 143520 240692 143540
rect 240692 143520 240744 143540
rect 240744 143520 240746 143540
rect 240874 143520 240930 143576
rect 240138 5072 240194 5128
rect 244186 240080 244242 240136
rect 244186 193160 244242 193216
rect 244186 173848 244242 173904
rect 244186 164212 244242 164248
rect 244186 164192 244188 164212
rect 244188 164192 244240 164212
rect 244240 164192 244242 164212
rect 244186 154536 244242 154592
rect 242898 5344 242954 5400
rect 242070 5208 242126 5264
rect 244370 258052 244426 258088
rect 244370 258032 244372 258052
rect 244372 258032 244424 258052
rect 244424 258032 244426 258052
rect 244370 240080 244426 240136
rect 244646 258032 244702 258088
rect 244462 193160 244518 193216
rect 244462 173884 244464 173904
rect 244464 173884 244516 173904
rect 244516 173884 244518 173904
rect 244462 173848 244518 173884
rect 244370 164212 244426 164248
rect 244370 164192 244372 164212
rect 244372 164192 244424 164212
rect 244424 164192 244426 164212
rect 244462 154536 244518 154592
rect 244462 138624 244518 138680
rect 244370 125568 244426 125624
rect 244922 164328 244978 164384
rect 245014 164192 245070 164248
rect 245842 183504 245898 183560
rect 245842 124208 245898 124264
rect 246026 183504 246082 183560
rect 246026 124208 246082 124264
rect 245750 5480 245806 5536
rect 246486 267824 246542 267880
rect 246762 267824 246818 267880
rect 246302 267688 246358 267744
rect 246486 267688 246542 267744
rect 246394 193196 246396 193216
rect 246396 193196 246448 193216
rect 246448 193196 246450 193216
rect 246394 193160 246450 193196
rect 246578 193196 246580 193216
rect 246580 193196 246632 193216
rect 246632 193196 246634 193216
rect 246578 193160 246634 193196
rect 246486 154672 246542 154728
rect 246394 154536 246450 154592
rect 246394 77560 246450 77616
rect 246394 77288 246450 77344
rect 246946 40432 247002 40488
rect 246946 40296 247002 40352
rect 249706 86964 249762 87000
rect 249706 86944 249708 86964
rect 249708 86944 249760 86964
rect 249760 86944 249762 86964
rect 252098 86808 252154 86864
rect 253018 269048 253074 269104
rect 253110 268912 253166 268968
rect 253018 230424 253074 230480
rect 253294 230424 253350 230480
rect 253018 211112 253074 211168
rect 253202 211112 253258 211168
rect 253110 26152 253166 26208
rect 253294 26152 253350 26208
rect 254490 29416 254546 29472
rect 254490 29008 254546 29064
rect 255042 328616 255098 328672
rect 254674 328480 254730 328536
rect 254766 164328 254822 164384
rect 254766 164192 254822 164248
rect 256698 328480 256754 328536
rect 257066 328480 257122 328536
rect 256974 124208 257030 124264
rect 257158 124208 257214 124264
rect 256606 40568 256662 40624
rect 256606 40160 256662 40216
rect 258814 298016 258870 298072
rect 258722 297880 258778 297936
rect 258630 230560 258686 230616
rect 258722 230424 258778 230480
rect 258814 164328 258870 164384
rect 258814 164192 258870 164248
rect 258722 93744 258778 93800
rect 258906 93744 258962 93800
rect 260194 248376 260250 248432
rect 260378 248376 260434 248432
rect 259458 86944 259514 87000
rect 259458 86808 259514 86864
rect 259458 40160 259514 40216
rect 259458 40024 259514 40080
rect 259458 17040 259514 17096
rect 259458 16632 259514 16688
rect 261390 278704 261446 278760
rect 261574 278704 261630 278760
rect 262954 336912 263010 336968
rect 262770 336776 262826 336832
rect 262862 200096 262918 200152
rect 263046 200096 263102 200152
rect 264334 269048 264390 269104
rect 264518 269084 264520 269104
rect 264520 269084 264572 269104
rect 264572 269084 264574 269104
rect 264518 269048 264574 269084
rect 264334 249736 264390 249792
rect 264518 249736 264574 249792
rect 264334 201476 264390 201512
rect 264334 201456 264336 201476
rect 264336 201456 264388 201476
rect 264388 201456 264390 201476
rect 264518 201476 264574 201512
rect 264518 201456 264520 201476
rect 264520 201456 264572 201476
rect 264572 201456 264574 201476
rect 264334 191820 264390 191856
rect 264334 191800 264336 191820
rect 264336 191800 264388 191820
rect 264388 191800 264390 191820
rect 264518 191820 264574 191856
rect 264518 191800 264520 191820
rect 264520 191800 264572 191820
rect 264572 191800 264574 191820
rect 264334 182144 264390 182200
rect 264518 182144 264574 182200
rect 264242 16224 264298 16280
rect 264242 15544 264298 15600
rect 266358 338136 266414 338192
rect 265622 269048 265678 269104
rect 265806 269084 265808 269104
rect 265808 269084 265860 269104
rect 265860 269084 265862 269104
rect 265806 269048 265862 269084
rect 265622 248376 265678 248432
rect 265806 248376 265862 248432
rect 265622 229064 265678 229120
rect 265806 229064 265862 229120
rect 265622 209752 265678 209808
rect 265806 209752 265862 209808
rect 265622 182144 265678 182200
rect 265806 182144 265862 182200
rect 265806 74568 265862 74624
rect 265622 64912 265678 64968
rect 265806 64912 265862 64968
rect 266910 328344 266966 328400
rect 266358 74568 266414 74624
rect 267554 5480 267610 5536
rect 267738 63552 267794 63608
rect 267738 63144 267794 63200
rect 267738 40432 267794 40488
rect 267738 40024 267794 40080
rect 268658 16360 268714 16416
rect 269026 16360 269082 16416
rect 268842 5072 268898 5128
rect 263414 3168 263470 3224
rect 263690 3168 263746 3224
rect 269026 5344 269082 5400
rect 270222 5208 270278 5264
rect 270406 4936 270462 4992
rect 270314 4800 270370 4856
rect 272246 336912 272302 336968
rect 272522 336776 272578 336832
rect 272338 336640 272394 336696
rect 272522 336640 272578 336696
rect 273074 4120 273130 4176
rect 273350 4120 273406 4176
rect 275190 3168 275246 3224
rect 278870 63688 278926 63744
rect 278962 63552 279018 63608
rect 278502 16496 278558 16552
rect 278686 16496 278742 16552
rect 278134 16224 278190 16280
rect 278686 16224 278742 16280
rect 282366 19216 282422 19272
rect 283562 40160 283618 40216
rect 283562 39752 283618 39808
rect 283562 19080 283618 19136
rect 284114 9560 284170 9616
rect 286690 19216 286746 19272
rect 287058 40160 287114 40216
rect 287058 39616 287114 39672
rect 288438 19080 288494 19136
rect 289358 13640 289414 13696
rect 289634 6704 289690 6760
rect 282826 3168 282882 3224
rect 290646 13504 290702 13560
rect 290830 13368 290886 13424
rect 291014 6568 291070 6624
rect 291934 13232 291990 13288
rect 292118 13096 292174 13152
rect 291106 6432 291162 6488
rect 292394 6296 292450 6352
rect 293130 288360 293186 288416
rect 293314 288396 293316 288416
rect 293316 288396 293368 288416
rect 293368 288396 293370 288416
rect 293314 288360 293370 288396
rect 293130 269048 293186 269104
rect 293314 269048 293370 269104
rect 293130 249736 293186 249792
rect 293314 249736 293370 249792
rect 293130 230424 293186 230480
rect 293314 230424 293370 230480
rect 293130 220804 293132 220824
rect 293132 220804 293184 220824
rect 293184 220804 293186 220824
rect 293130 220768 293186 220804
rect 293314 220804 293316 220824
rect 293316 220804 293368 220824
rect 293368 220804 293370 220824
rect 293314 220768 293370 220804
rect 293130 211132 293186 211168
rect 293130 211112 293132 211132
rect 293132 211112 293184 211132
rect 293184 211112 293186 211132
rect 293314 211132 293370 211168
rect 293314 211112 293316 211132
rect 293316 211112 293368 211132
rect 293368 211112 293370 211132
rect 293130 201476 293186 201512
rect 293130 201456 293132 201476
rect 293132 201456 293184 201476
rect 293184 201456 293186 201476
rect 293314 201476 293370 201512
rect 293314 201456 293316 201476
rect 293316 201456 293368 201476
rect 293368 201456 293370 201476
rect 293130 191820 293186 191856
rect 293130 191800 293132 191820
rect 293132 191800 293184 191820
rect 293184 191800 293186 191820
rect 293314 191820 293370 191856
rect 293314 191800 293316 191820
rect 293316 191800 293368 191820
rect 293368 191800 293370 191820
rect 293130 182164 293186 182200
rect 293130 182144 293132 182164
rect 293132 182144 293184 182164
rect 293184 182144 293186 182164
rect 293314 182164 293370 182200
rect 293314 182144 293316 182164
rect 293316 182144 293368 182164
rect 293368 182144 293370 182164
rect 292578 17040 292634 17096
rect 292578 16768 292634 16824
rect 294786 211248 294842 211304
rect 294786 211132 294842 211168
rect 294786 211112 294788 211132
rect 294788 211112 294840 211132
rect 294840 211112 294842 211132
rect 294602 201456 294658 201512
rect 294786 201456 294842 201512
rect 294786 191936 294842 191992
rect 294786 191820 294842 191856
rect 294786 191800 294788 191820
rect 294788 191800 294840 191820
rect 294840 191800 294842 191820
rect 294602 182144 294658 182200
rect 294786 182144 294842 182200
rect 296074 211248 296130 211304
rect 296074 211132 296130 211168
rect 296074 211112 296076 211132
rect 296076 211112 296128 211132
rect 296128 211112 296130 211132
rect 295890 201456 295946 201512
rect 296074 201456 296130 201512
rect 296074 191936 296130 191992
rect 296074 191820 296130 191856
rect 296074 191800 296076 191820
rect 296076 191800 296128 191820
rect 296128 191800 296130 191820
rect 295890 182144 295946 182200
rect 296074 182144 296130 182200
rect 292486 6160 292542 6216
rect 292394 4120 292450 4176
rect 292670 4120 292726 4176
rect 297362 16224 297418 16280
rect 297362 15544 297418 15600
rect 300490 10784 300546 10840
rect 300582 10648 300638 10704
rect 301594 218048 301650 218104
rect 301778 218048 301834 218104
rect 301594 198736 301650 198792
rect 301778 198736 301834 198792
rect 301962 141208 302018 141264
rect 301962 140800 302018 140856
rect 300858 17040 300914 17096
rect 300858 16904 300914 16960
rect 301962 10512 302018 10568
rect 303434 10376 303490 10432
rect 303342 10240 303398 10296
rect 305182 336912 305238 336968
rect 305366 336776 305422 336832
rect 305918 17720 305974 17776
rect 308402 16224 308458 16280
rect 308402 15544 308458 15600
rect 308770 8200 308826 8256
rect 310242 8064 310298 8120
rect 310150 7928 310206 7984
rect 309782 5480 309838 5536
rect 311530 7792 311586 7848
rect 311990 16768 312046 16824
rect 311898 16632 311954 16688
rect 312910 7656 312966 7712
rect 313002 7520 313058 7576
rect 314198 17584 314254 17640
rect 313370 5344 313426 5400
rect 311806 4120 311862 4176
rect 315578 17448 315634 17504
rect 315486 17312 315542 17368
rect 313922 4120 313978 4176
rect 315762 5072 315818 5128
rect 318154 335280 318210 335336
rect 318430 335280 318486 335336
rect 317142 9424 317198 9480
rect 317050 5208 317106 5264
rect 318430 9288 318486 9344
rect 319442 325660 319444 325680
rect 319444 325660 319496 325680
rect 319496 325660 319498 325680
rect 319442 325624 319498 325660
rect 319626 325624 319682 325680
rect 319442 277344 319498 277400
rect 319626 277344 319682 277400
rect 319442 229064 319498 229120
rect 319626 229064 319682 229120
rect 319626 143656 319682 143712
rect 319626 143520 319682 143576
rect 319718 12280 319774 12336
rect 319534 12144 319590 12200
rect 319810 9152 319866 9208
rect 319902 9016 319958 9072
rect 319994 5480 320050 5536
rect 319258 4936 319314 4992
rect 320914 278704 320970 278760
rect 321098 278704 321154 278760
rect 320914 269084 320916 269104
rect 320916 269084 320968 269104
rect 320968 269084 320970 269104
rect 320914 269048 320970 269084
rect 321098 269084 321100 269104
rect 321100 269084 321152 269104
rect 321152 269084 321154 269104
rect 321098 269048 321154 269084
rect 320914 259428 320916 259448
rect 320916 259428 320968 259448
rect 320968 259428 320970 259448
rect 320914 259392 320970 259428
rect 321098 259428 321100 259448
rect 321100 259428 321152 259448
rect 321152 259428 321154 259448
rect 321098 259392 321154 259428
rect 320914 249772 320916 249792
rect 320916 249772 320968 249792
rect 320968 249772 320970 249792
rect 320914 249736 320970 249772
rect 321098 249772 321100 249792
rect 321100 249772 321152 249792
rect 321152 249772 321154 249792
rect 321098 249736 321154 249772
rect 320914 240116 320916 240136
rect 320916 240116 320968 240136
rect 320968 240116 320970 240136
rect 320914 240080 320970 240116
rect 321098 240116 321100 240136
rect 321100 240116 321152 240136
rect 321152 240116 321154 240136
rect 321098 240080 321154 240116
rect 320914 230460 320916 230480
rect 320916 230460 320968 230480
rect 320968 230460 320970 230480
rect 320914 230424 320970 230460
rect 321098 230460 321100 230480
rect 321100 230460 321152 230480
rect 321152 230460 321154 230480
rect 321098 230424 321154 230460
rect 321098 201592 321154 201648
rect 321098 201456 321154 201512
rect 321098 182280 321154 182336
rect 321098 182144 321154 182200
rect 320914 142160 320970 142216
rect 321006 141888 321062 141944
rect 320914 113192 320970 113248
rect 321098 113192 321154 113248
rect 321006 12008 321062 12064
rect 321190 8880 321246 8936
rect 321282 6840 321338 6896
rect 321374 5344 321430 5400
rect 322018 337184 322074 337240
rect 322294 259428 322296 259448
rect 322296 259428 322348 259448
rect 322348 259428 322350 259448
rect 322294 259392 322350 259428
rect 322202 259256 322258 259312
rect 322110 248376 322166 248432
rect 322294 248376 322350 248432
rect 322110 229064 322166 229120
rect 322294 229064 322350 229120
rect 322110 219408 322166 219464
rect 322294 219408 322350 219464
rect 322110 201456 322166 201512
rect 322294 201456 322350 201512
rect 322294 161336 322350 161392
rect 322386 161200 322442 161256
rect 322294 11872 322350 11928
rect 322478 11192 322534 11248
rect 321466 5208 321522 5264
rect 322662 5072 322718 5128
rect 322938 16768 322994 16824
rect 323306 11736 323362 11792
rect 323950 337184 324006 337240
rect 323950 11736 324006 11792
rect 323398 11600 323454 11656
rect 324042 11600 324098 11656
rect 322846 4936 322902 4992
rect 322846 4800 322902 4856
rect 324226 4800 324282 4856
rect 324594 15816 324650 15872
rect 326158 337456 326214 337512
rect 325974 337320 326030 337376
rect 325882 16088 325938 16144
rect 325790 14592 325846 14648
rect 324778 14456 324834 14512
rect 324410 12960 324466 13016
rect 324318 3304 324374 3360
rect 324870 4120 324926 4176
rect 326250 296656 326306 296712
rect 326434 296656 326490 296712
rect 326250 277344 326306 277400
rect 326526 277344 326582 277400
rect 326158 15952 326214 16008
rect 327078 6840 327134 6896
rect 326066 3440 326122 3496
rect 327354 16360 327410 16416
rect 327446 16224 327502 16280
rect 327262 3712 327318 3768
rect 327538 3576 327594 3632
rect 328182 337592 328238 337648
rect 328642 10920 328698 10976
rect 328550 3984 328606 4040
rect 329010 298016 329066 298072
rect 329194 298016 329250 298072
rect 329010 288360 329066 288416
rect 329194 288360 329250 288416
rect 329010 62056 329066 62112
rect 329194 62056 329250 62112
rect 329194 34448 329250 34504
rect 329378 34448 329434 34504
rect 328826 17992 328882 18048
rect 328734 3848 328790 3904
rect 331310 337728 331366 337784
rect 330758 335280 330814 335336
rect 330942 335280 330998 335336
rect 330574 247288 330630 247344
rect 330574 247036 330630 247072
rect 330574 247016 330576 247036
rect 330576 247016 330628 247036
rect 330628 247016 330630 247036
rect 330758 215328 330814 215384
rect 330942 215328 330998 215384
rect 330758 205672 330814 205728
rect 330942 205672 330998 205728
rect 331586 256672 331642 256728
rect 330298 4120 330354 4176
rect 331770 256672 331826 256728
rect 331770 237360 331826 237416
rect 331954 237360 332010 237416
rect 332506 16904 332562 16960
rect 333242 247152 333298 247208
rect 333242 247036 333298 247072
rect 333242 247016 333244 247036
rect 333244 247016 333296 247036
rect 333296 247016 333298 247036
rect 333242 237360 333298 237416
rect 333426 237360 333482 237416
rect 333886 63960 333942 64016
rect 333886 63688 333942 63744
rect 333886 40296 333942 40352
rect 333886 40160 333942 40216
rect 333886 16904 333942 16960
rect 333886 16632 333942 16688
rect 334162 14864 334218 14920
rect 333242 14728 333298 14784
rect 335450 40160 335506 40216
rect 334530 15000 334586 15056
rect 335818 288360 335874 288416
rect 336002 288360 336058 288416
rect 335818 238720 335874 238776
rect 336002 238720 336058 238776
rect 335910 190440 335966 190496
rect 336094 190440 336150 190496
rect 335910 161472 335966 161528
rect 336094 161472 336150 161528
rect 335634 15136 335690 15192
rect 337934 29280 337990 29336
rect 338118 29280 338174 29336
rect 338394 17176 338450 17232
rect 340050 270680 340106 270736
rect 340326 270408 340382 270464
rect 339958 230460 339960 230480
rect 339960 230460 340012 230480
rect 340012 230460 340014 230480
rect 339958 230424 340014 230460
rect 340142 230424 340198 230480
rect 340142 164212 340198 164248
rect 340142 164192 340144 164212
rect 340144 164192 340196 164212
rect 340196 164192 340198 164212
rect 340326 164192 340382 164248
rect 340142 144880 340198 144936
rect 340418 144880 340474 144936
rect 341706 211112 341762 211168
rect 341890 211112 341946 211168
rect 344926 40316 344982 40352
rect 344926 40296 344928 40316
rect 344928 40296 344980 40316
rect 344980 40296 344982 40316
rect 345018 16244 345074 16280
rect 345018 16224 345020 16244
rect 345020 16224 345072 16244
rect 345072 16224 345074 16244
rect 345386 259392 345442 259448
rect 345570 259392 345626 259448
rect 345386 191800 345442 191856
rect 345570 191800 345626 191856
rect 345386 154536 345442 154592
rect 345570 154536 345626 154592
rect 345294 124208 345350 124264
rect 345570 124208 345626 124264
rect 346398 16496 346454 16552
rect 371882 310936 371938 310992
rect 350446 310664 350502 310720
rect 367006 310664 367062 310720
rect 350630 310528 350686 310584
rect 371882 310528 371938 310584
rect 367006 310256 367062 310312
rect 371882 264016 371938 264072
rect 350446 263744 350502 263800
rect 367006 263744 367062 263800
rect 350630 263608 350686 263664
rect 371882 263608 371938 263664
rect 367006 263336 367062 263392
rect 371882 217096 371938 217152
rect 350446 216824 350502 216880
rect 367006 216824 367062 216880
rect 350630 216688 350686 216744
rect 371882 216688 371938 216744
rect 367006 216416 367062 216472
rect 371882 170176 371938 170232
rect 350446 169904 350502 169960
rect 367006 169904 367062 169960
rect 350630 169768 350686 169824
rect 371882 169768 371938 169824
rect 367006 169496 367062 169552
rect 579802 457816 579858 457872
rect 579802 439864 579858 439920
rect 579802 404776 579858 404832
rect 579894 357856 579950 357912
rect 579986 322632 580042 322688
rect 580170 451696 580226 451752
rect 580078 299104 580134 299160
rect 580170 275712 580226 275768
rect 579618 123120 579674 123176
rect 375286 87352 375342 87408
rect 350446 87080 350502 87136
rect 360290 87080 360346 87136
rect 350630 86944 350686 87000
rect 360106 86944 360162 87000
rect 386326 87216 386382 87272
rect 379426 87116 379428 87136
rect 379428 87116 379480 87136
rect 379480 87116 379482 87136
rect 379426 87080 379482 87116
rect 375286 86944 375342 87000
rect 580906 252184 580962 252240
rect 580814 228792 580870 228848
rect 580722 205264 580778 205320
rect 580630 181872 580686 181928
rect 580538 158344 580594 158400
rect 580446 134816 580502 134872
rect 580354 111424 580410 111480
rect 580262 76200 580318 76256
rect 353206 63960 353262 64016
rect 371882 63960 371938 64016
rect 353206 63688 353262 63744
rect 354586 63688 354642 63744
rect 367006 63688 367062 63744
rect 354586 63552 354642 63608
rect 364246 63416 364302 63472
rect 371882 63552 371938 63608
rect 364246 63280 364302 63336
rect 367006 63280 367062 63336
rect 355966 40568 356022 40624
rect 371882 40432 371938 40488
rect 367006 40160 367062 40216
rect 355966 40024 356022 40080
rect 371882 40024 371938 40080
rect 367006 39752 367062 39808
rect 355966 29416 356022 29472
rect 375286 29416 375342 29472
rect 360290 29144 360346 29200
rect 386326 29280 386382 29336
rect 379426 29180 379428 29200
rect 379428 29180 379480 29200
rect 379480 29180 379482 29200
rect 379426 29144 379482 29180
rect 355966 29008 356022 29064
rect 360106 29008 360162 29064
rect 375286 29008 375342 29064
rect 369766 16768 369822 16824
rect 379610 16768 379666 16824
rect 369950 16632 370006 16688
rect 379426 16632 379482 16688
rect 384670 9560 384726 9616
rect 389086 16768 389142 16824
rect 389270 16632 389326 16688
rect 404266 16768 404322 16824
rect 408406 16768 408462 16824
rect 394698 16668 394700 16688
rect 394700 16668 394752 16688
rect 394752 16668 394754 16688
rect 394698 16632 394754 16668
rect 408590 16632 408646 16688
rect 414018 13640 414074 13696
rect 416778 13504 416834 13560
rect 415674 6704 415730 6760
rect 420918 13368 420974 13424
rect 419170 6568 419226 6624
rect 425058 13232 425114 13288
rect 422758 6432 422814 6488
rect 427818 13096 427874 13152
rect 426346 6296 426402 6352
rect 429934 6160 429990 6216
rect 437386 16652 437442 16688
rect 437386 16632 437388 16652
rect 437388 16632 437440 16652
rect 437440 16632 437442 16652
rect 442906 16652 442962 16688
rect 442906 16632 442908 16652
rect 442908 16632 442960 16652
rect 442960 16632 442962 16652
rect 492678 17720 492734 17776
rect 447046 16768 447102 16824
rect 447230 16768 447286 16824
rect 466366 16768 466422 16824
rect 476210 16768 476266 16824
rect 466550 16632 466606 16688
rect 476026 16632 476082 16688
rect 466458 10784 466514 10840
rect 469218 10648 469274 10704
rect 473358 10512 473414 10568
rect 477590 10376 477646 10432
rect 480258 10240 480314 10296
rect 491206 16768 491262 16824
rect 491206 16496 491262 16552
rect 534078 17584 534134 17640
rect 495346 17040 495402 17096
rect 495530 17040 495586 17096
rect 505006 16924 505062 16960
rect 505006 16904 505008 16924
rect 505008 16904 505060 16924
rect 505060 16904 505062 16924
rect 511906 16768 511962 16824
rect 509606 8200 509662 8256
rect 513194 8064 513250 8120
rect 516782 7928 516838 7984
rect 523866 7792 523922 7848
rect 527454 7656 527510 7712
rect 531042 7520 531098 7576
rect 536838 17448 536894 17504
rect 540978 17312 541034 17368
rect 560298 12280 560354 12336
rect 548890 9424 548946 9480
rect 555974 9288 556030 9344
rect 559562 9152 559618 9208
rect 563058 12144 563114 12200
rect 561954 5480 562010 5536
rect 567198 12008 567254 12064
rect 563150 9016 563206 9072
rect 565542 5344 565598 5400
rect 574098 11872 574154 11928
rect 570234 8880 570290 8936
rect 569038 5208 569094 5264
rect 572626 5072 572682 5128
rect 578238 11736 578294 11792
rect 576214 4936 576270 4992
rect 580998 11600 581054 11656
rect 579802 4800 579858 4856
<< metal3 >>
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect 494881 686082 494947 686085
rect 494102 686080 494947 686082
rect 494102 686024 494886 686080
rect 494942 686024 494947 686080
rect 494102 686022 494947 686024
rect 494102 685946 494162 686022
rect 494881 686019 494947 686022
rect 494237 685946 494303 685949
rect 494102 685944 494303 685946
rect 494102 685888 494242 685944
rect 494298 685888 494303 685944
rect 494102 685886 494303 685888
rect 494237 685883 494303 685886
rect -960 682274 480 682364
rect 3509 682274 3575 682277
rect -960 682272 3575 682274
rect -960 682216 3514 682272
rect 3570 682216 3575 682272
rect -960 682214 3575 682216
rect -960 682124 480 682214
rect 3509 682211 3575 682214
rect 580165 674658 580231 674661
rect 583520 674658 584960 674748
rect 580165 674656 584960 674658
rect 580165 674600 580170 674656
rect 580226 674600 584960 674656
rect 580165 674598 584960 674600
rect 580165 674595 580231 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 580165 651130 580231 651133
rect 583520 651130 584960 651220
rect 580165 651128 584960 651130
rect 580165 651072 580170 651128
rect 580226 651072 584960 651128
rect 580165 651070 584960 651072
rect 580165 651067 580231 651070
rect 583520 650980 584960 651070
rect 580165 639434 580231 639437
rect 583520 639434 584960 639524
rect 580165 639432 584960 639434
rect 580165 639376 580170 639432
rect 580226 639376 584960 639432
rect 580165 639374 584960 639376
rect 580165 639371 580231 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 580165 627738 580231 627741
rect 583520 627738 584960 627828
rect 580165 627736 584960 627738
rect 580165 627680 580170 627736
rect 580226 627680 584960 627736
rect 580165 627678 584960 627680
rect 580165 627675 580231 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3417 624882 3483 624885
rect -960 624880 3483 624882
rect -960 624824 3422 624880
rect 3478 624824 3483 624880
rect -960 624822 3483 624824
rect -960 624732 480 624822
rect 3417 624819 3483 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3417 610466 3483 610469
rect -960 610464 3483 610466
rect -960 610408 3422 610464
rect 3478 610408 3483 610464
rect -960 610406 3483 610408
rect -960 610316 480 610406
rect 3417 610403 3483 610406
rect 580165 604210 580231 604213
rect 583520 604210 584960 604300
rect 580165 604208 584960 604210
rect 580165 604152 580170 604208
rect 580226 604152 584960 604208
rect 580165 604150 584960 604152
rect 580165 604147 580231 604150
rect 583520 604060 584960 604150
rect -960 596050 480 596140
rect 3233 596050 3299 596053
rect -960 596048 3299 596050
rect -960 595992 3238 596048
rect 3294 595992 3299 596048
rect -960 595990 3299 595992
rect -960 595900 480 595990
rect 3233 595987 3299 595990
rect 580165 592514 580231 592517
rect 583520 592514 584960 592604
rect 580165 592512 584960 592514
rect 580165 592456 580170 592512
rect 580226 592456 584960 592512
rect 580165 592454 584960 592456
rect 580165 592451 580231 592454
rect 583520 592364 584960 592454
rect -960 581620 480 581860
rect 580165 580818 580231 580821
rect 583520 580818 584960 580908
rect 580165 580816 584960 580818
rect 580165 580760 580170 580816
rect 580226 580760 584960 580816
rect 580165 580758 584960 580760
rect 580165 580755 580231 580758
rect 583520 580668 584960 580758
rect 493869 579730 493935 579733
rect 494053 579730 494119 579733
rect 493869 579728 494119 579730
rect 493869 579672 493874 579728
rect 493930 579672 494058 579728
rect 494114 579672 494119 579728
rect 493869 579670 494119 579672
rect 493869 579667 493935 579670
rect 494053 579667 494119 579670
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3417 567354 3483 567357
rect -960 567352 3483 567354
rect -960 567296 3422 567352
rect 3478 567296 3483 567352
rect -960 567294 3483 567296
rect -960 567204 480 567294
rect 3417 567291 3483 567294
rect 494145 560282 494211 560285
rect 494329 560282 494395 560285
rect 494145 560280 494395 560282
rect 494145 560224 494150 560280
rect 494206 560224 494334 560280
rect 494390 560224 494395 560280
rect 494145 560222 494395 560224
rect 494145 560219 494211 560222
rect 494329 560219 494395 560222
rect 580165 557290 580231 557293
rect 583520 557290 584960 557380
rect 580165 557288 584960 557290
rect 580165 557232 580170 557288
rect 580226 557232 584960 557288
rect 580165 557230 584960 557232
rect 580165 557227 580231 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 3141 553074 3207 553077
rect -960 553072 3207 553074
rect -960 553016 3146 553072
rect 3202 553016 3207 553072
rect -960 553014 3207 553016
rect -960 552924 480 553014
rect 3141 553011 3207 553014
rect 580165 545594 580231 545597
rect 583520 545594 584960 545684
rect 580165 545592 584960 545594
rect 580165 545536 580170 545592
rect 580226 545536 584960 545592
rect 580165 545534 584960 545536
rect 580165 545531 580231 545534
rect 583520 545444 584960 545534
rect 218973 540970 219039 540973
rect 219157 540970 219223 540973
rect 218973 540968 219223 540970
rect 218973 540912 218978 540968
rect 219034 540912 219162 540968
rect 219218 540912 219223 540968
rect 218973 540910 219223 540912
rect 218973 540907 219039 540910
rect 219157 540907 219223 540910
rect 494145 540970 494211 540973
rect 494329 540970 494395 540973
rect 494145 540968 494395 540970
rect 494145 540912 494150 540968
rect 494206 540912 494334 540968
rect 494390 540912 494395 540968
rect 494145 540910 494395 540912
rect 494145 540907 494211 540910
rect 494329 540907 494395 540910
rect -960 538658 480 538748
rect 3417 538658 3483 538661
rect -960 538656 3483 538658
rect -960 538600 3422 538656
rect 3478 538600 3483 538656
rect -960 538598 3483 538600
rect -960 538508 480 538598
rect 3417 538595 3483 538598
rect 580165 533898 580231 533901
rect 583520 533898 584960 533988
rect 580165 533896 584960 533898
rect 580165 533840 580170 533896
rect 580226 533840 584960 533896
rect 580165 533838 584960 533840
rect 580165 533835 580231 533838
rect 583520 533748 584960 533838
rect 218973 531314 219039 531317
rect 219157 531314 219223 531317
rect 218973 531312 219223 531314
rect 218973 531256 218978 531312
rect 219034 531256 219162 531312
rect 219218 531256 219223 531312
rect 218973 531254 219223 531256
rect 218973 531251 219039 531254
rect 219157 531251 219223 531254
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 218789 521658 218855 521661
rect 218973 521658 219039 521661
rect 218789 521656 219039 521658
rect 218789 521600 218794 521656
rect 218850 521600 218978 521656
rect 219034 521600 219039 521656
rect 218789 521598 219039 521600
rect 218789 521595 218855 521598
rect 218973 521595 219039 521598
rect 494145 521658 494211 521661
rect 494329 521658 494395 521661
rect 494145 521656 494395 521658
rect 494145 521600 494150 521656
rect 494206 521600 494334 521656
rect 494390 521600 494395 521656
rect 494145 521598 494395 521600
rect 494145 521595 494211 521598
rect 494329 521595 494395 521598
rect 542537 521658 542603 521661
rect 542721 521658 542787 521661
rect 542537 521656 542787 521658
rect 542537 521600 542542 521656
rect 542598 521600 542726 521656
rect 542782 521600 542787 521656
rect 542537 521598 542787 521600
rect 542537 521595 542603 521598
rect 542721 521595 542787 521598
rect 559097 521658 559163 521661
rect 559281 521658 559347 521661
rect 559097 521656 559347 521658
rect 559097 521600 559102 521656
rect 559158 521600 559286 521656
rect 559342 521600 559347 521656
rect 559097 521598 559347 521600
rect 559097 521595 559163 521598
rect 559281 521595 559347 521598
rect 580165 510370 580231 510373
rect 583520 510370 584960 510460
rect 580165 510368 584960 510370
rect 580165 510312 580170 510368
rect 580226 510312 584960 510368
rect 580165 510310 584960 510312
rect 580165 510307 580231 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3417 509962 3483 509965
rect -960 509960 3483 509962
rect -960 509904 3422 509960
rect 3478 509904 3483 509960
rect -960 509902 3483 509904
rect -960 509812 480 509902
rect 3417 509899 3483 509902
rect 493961 502346 494027 502349
rect 494237 502346 494303 502349
rect 493961 502344 494303 502346
rect 493961 502288 493966 502344
rect 494022 502288 494242 502344
rect 494298 502288 494303 502344
rect 493961 502286 494303 502288
rect 493961 502283 494027 502286
rect 494237 502283 494303 502286
rect 542353 502346 542419 502349
rect 542629 502346 542695 502349
rect 542353 502344 542695 502346
rect 542353 502288 542358 502344
rect 542414 502288 542634 502344
rect 542690 502288 542695 502344
rect 542353 502286 542695 502288
rect 542353 502283 542419 502286
rect 542629 502283 542695 502286
rect 558913 502346 558979 502349
rect 559189 502346 559255 502349
rect 558913 502344 559255 502346
rect 558913 502288 558918 502344
rect 558974 502288 559194 502344
rect 559250 502288 559255 502344
rect 558913 502286 559255 502288
rect 558913 502283 558979 502286
rect 559189 502283 559255 502286
rect 580165 498674 580231 498677
rect 583520 498674 584960 498764
rect 580165 498672 584960 498674
rect 580165 498616 580170 498672
rect 580226 498616 584960 498672
rect 580165 498614 584960 498616
rect 580165 498611 580231 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 3417 495546 3483 495549
rect -960 495544 3483 495546
rect -960 495488 3422 495544
rect 3478 495488 3483 495544
rect -960 495486 3483 495488
rect -960 495396 480 495486
rect 3417 495483 3483 495486
rect 493961 492690 494027 492693
rect 494145 492690 494211 492693
rect 493961 492688 494211 492690
rect 493961 492632 493966 492688
rect 494022 492632 494150 492688
rect 494206 492632 494211 492688
rect 493961 492630 494211 492632
rect 493961 492627 494027 492630
rect 494145 492627 494211 492630
rect 542353 492690 542419 492693
rect 542537 492690 542603 492693
rect 542353 492688 542603 492690
rect 542353 492632 542358 492688
rect 542414 492632 542542 492688
rect 542598 492632 542603 492688
rect 542353 492630 542603 492632
rect 542353 492627 542419 492630
rect 542537 492627 542603 492630
rect 558913 492690 558979 492693
rect 559097 492690 559163 492693
rect 558913 492688 559163 492690
rect 558913 492632 558918 492688
rect 558974 492632 559102 492688
rect 559158 492632 559163 492688
rect 558913 492630 559163 492632
rect 558913 492627 558979 492630
rect 559097 492627 559163 492630
rect 580165 486842 580231 486845
rect 583520 486842 584960 486932
rect 580165 486840 584960 486842
rect 580165 486784 580170 486840
rect 580226 486784 584960 486840
rect 580165 486782 584960 486784
rect 580165 486779 580231 486782
rect 583520 486692 584960 486782
rect -960 481130 480 481220
rect 3141 481130 3207 481133
rect -960 481128 3207 481130
rect -960 481072 3146 481128
rect 3202 481072 3207 481128
rect -960 481070 3207 481072
rect -960 480980 480 481070
rect 3141 481067 3207 481070
rect 583520 474996 584960 475236
rect -960 466700 480 466940
rect 154297 463722 154363 463725
rect 154481 463722 154547 463725
rect 154297 463720 154547 463722
rect 154297 463664 154302 463720
rect 154358 463664 154486 463720
rect 154542 463664 154547 463720
rect 154297 463662 154547 463664
rect 154297 463659 154363 463662
rect 154481 463659 154547 463662
rect 580073 463450 580139 463453
rect 583520 463450 584960 463540
rect 580073 463448 584960 463450
rect 580073 463392 580078 463448
rect 580134 463392 584960 463448
rect 580073 463390 584960 463392
rect 580073 463387 580139 463390
rect 583520 463300 584960 463390
rect 252461 463042 252527 463045
rect 348366 463042 348372 463044
rect 252461 463040 348372 463042
rect 252461 462984 252466 463040
rect 252522 462984 348372 463040
rect 252461 462982 348372 462984
rect 252461 462979 252527 462982
rect 348366 462980 348372 462982
rect 348436 462980 348442 463044
rect 232446 462844 232452 462908
rect 232516 462906 232522 462908
rect 318701 462906 318767 462909
rect 232516 462904 318767 462906
rect 232516 462848 318706 462904
rect 318762 462848 318767 462904
rect 232516 462846 318767 462848
rect 232516 462844 232522 462846
rect 318701 462843 318767 462846
rect 255589 462770 255655 462773
rect 348734 462770 348740 462772
rect 255589 462768 348740 462770
rect 255589 462712 255594 462768
rect 255650 462712 348740 462768
rect 255589 462710 348740 462712
rect 255589 462707 255655 462710
rect 348734 462708 348740 462710
rect 348804 462708 348810 462772
rect 256601 462634 256667 462637
rect 348918 462634 348924 462636
rect 256601 462632 348924 462634
rect 256601 462576 256606 462632
rect 256662 462576 348924 462632
rect 256601 462574 348924 462576
rect 256601 462571 256667 462574
rect 348918 462572 348924 462574
rect 348988 462572 348994 462636
rect 253473 462498 253539 462501
rect 348550 462498 348556 462500
rect 253473 462496 348556 462498
rect 253473 462440 253478 462496
rect 253534 462440 348556 462496
rect 253473 462438 348556 462440
rect 253473 462435 253539 462438
rect 348550 462436 348556 462438
rect 348620 462436 348626 462500
rect 251633 460050 251699 460053
rect 344318 460050 344324 460052
rect 251633 460048 344324 460050
rect 251633 459992 251638 460048
rect 251694 459992 344324 460048
rect 251633 459990 344324 459992
rect 251633 459987 251699 459990
rect 344318 459988 344324 459990
rect 344388 459988 344394 460052
rect 248321 459914 248387 459917
rect 344134 459914 344140 459916
rect 248321 459912 344140 459914
rect 248321 459856 248326 459912
rect 248382 459856 344140 459912
rect 248321 459854 344140 459856
rect 248321 459851 248387 459854
rect 344134 459852 344140 459854
rect 344204 459852 344210 459916
rect 245377 459778 245443 459781
rect 342478 459778 342484 459780
rect 245377 459776 342484 459778
rect 245377 459720 245382 459776
rect 245438 459720 342484 459776
rect 245377 459718 342484 459720
rect 245377 459715 245443 459718
rect 342478 459716 342484 459718
rect 342548 459716 342554 459780
rect 231669 459644 231735 459645
rect 231669 459640 231716 459644
rect 231780 459642 231786 459644
rect 232681 459642 232747 459645
rect 232998 459642 233004 459644
rect 231669 459584 231674 459640
rect 231669 459580 231716 459584
rect 231780 459582 231826 459642
rect 232681 459640 233004 459642
rect 232681 459584 232686 459640
rect 232742 459584 233004 459640
rect 232681 459582 233004 459584
rect 231780 459580 231786 459582
rect 231669 459579 231735 459580
rect 232681 459579 232747 459582
rect 232998 459580 233004 459582
rect 233068 459580 233074 459644
rect 233785 459642 233851 459645
rect 233918 459642 233924 459644
rect 233785 459640 233924 459642
rect 233785 459584 233790 459640
rect 233846 459584 233924 459640
rect 233785 459582 233924 459584
rect 233785 459579 233851 459582
rect 233918 459580 233924 459582
rect 233988 459580 233994 459644
rect 242249 459642 242315 459645
rect 342662 459642 342668 459644
rect 242249 459640 342668 459642
rect 242249 459584 242254 459640
rect 242310 459584 342668 459640
rect 242249 459582 342668 459584
rect 242249 459579 242315 459582
rect 342662 459580 342668 459582
rect 342732 459580 342738 459644
rect 343582 459580 343588 459644
rect 343652 459642 343658 459644
rect 343725 459642 343791 459645
rect 343652 459640 343791 459642
rect 343652 459584 343730 459640
rect 343786 459584 343791 459640
rect 343652 459582 343791 459584
rect 343652 459580 343658 459582
rect 343725 459579 343791 459582
rect 345289 459642 345355 459645
rect 345422 459642 345428 459644
rect 345289 459640 345428 459642
rect 345289 459584 345294 459640
rect 345350 459584 345428 459640
rect 345289 459582 345428 459584
rect 345289 459579 345355 459582
rect 345422 459580 345428 459582
rect 345492 459580 345498 459644
rect 233734 459308 233740 459372
rect 233804 459370 233810 459372
rect 234337 459370 234403 459373
rect 233804 459368 234403 459370
rect 233804 459312 234342 459368
rect 234398 459312 234403 459368
rect 233804 459310 234403 459312
rect 233804 459308 233810 459310
rect 234337 459307 234403 459310
rect 258809 459370 258875 459373
rect 258942 459370 258948 459372
rect 258809 459368 258948 459370
rect 258809 459312 258814 459368
rect 258870 459312 258948 459368
rect 258809 459310 258948 459312
rect 258809 459307 258875 459310
rect 258942 459308 258948 459310
rect 259012 459308 259018 459372
rect 324630 459308 324636 459372
rect 324700 459370 324706 459372
rect 324865 459370 324931 459373
rect 324700 459368 324931 459370
rect 324700 459312 324870 459368
rect 324926 459312 324931 459368
rect 324700 459310 324931 459312
rect 324700 459308 324706 459310
rect 324865 459307 324931 459310
rect 345238 459308 345244 459372
rect 345308 459370 345314 459372
rect 345749 459370 345815 459373
rect 345308 459368 345815 459370
rect 345308 459312 345754 459368
rect 345810 459312 345815 459368
rect 345308 459310 345815 459312
rect 345308 459308 345314 459310
rect 345749 459307 345815 459310
rect 347078 459308 347084 459372
rect 347148 459370 347154 459372
rect 347221 459370 347287 459373
rect 347148 459368 347287 459370
rect 347148 459312 347226 459368
rect 347282 459312 347287 459368
rect 347148 459310 347287 459312
rect 347148 459308 347154 459310
rect 347221 459307 347287 459310
rect 258942 457812 258948 457876
rect 259012 457874 259018 457876
rect 579797 457874 579863 457877
rect 259012 457872 579863 457874
rect 259012 457816 579802 457872
rect 579858 457816 579863 457872
rect 259012 457814 579863 457816
rect 259012 457812 259018 457814
rect 579797 457811 579863 457814
rect 3325 457738 3391 457741
rect 324630 457738 324636 457740
rect 3325 457736 324636 457738
rect 3325 457680 3330 457736
rect 3386 457680 324636 457736
rect 3325 457678 324636 457680
rect 3325 457675 3391 457678
rect 324630 457676 324636 457678
rect 324700 457676 324706 457740
rect 232446 452570 232452 452572
rect -960 452434 480 452524
rect 614 452510 232452 452570
rect 614 452434 674 452510
rect 232446 452508 232452 452510
rect 232516 452508 232522 452572
rect -960 452374 674 452434
rect -960 452284 480 452374
rect 580165 451754 580231 451757
rect 583520 451754 584960 451844
rect 580165 451752 584960 451754
rect 580165 451696 580170 451752
rect 580226 451696 584960 451752
rect 580165 451694 584960 451696
rect 580165 451691 580231 451694
rect 583520 451604 584960 451694
rect 579797 439922 579863 439925
rect 583520 439922 584960 440012
rect 579797 439920 584960 439922
rect 579797 439864 579802 439920
rect 579858 439864 584960 439920
rect 579797 439862 584960 439864
rect 579797 439859 579863 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 2773 438018 2839 438021
rect -960 438016 2839 438018
rect -960 437960 2778 438016
rect 2834 437960 2839 438016
rect -960 437958 2839 437960
rect -960 437868 480 437958
rect 2773 437955 2839 437958
rect 583520 428076 584960 428316
rect -960 423738 480 423828
rect 2957 423738 3023 423741
rect -960 423736 3023 423738
rect -960 423680 2962 423736
rect 3018 423680 3023 423736
rect -960 423678 3023 423680
rect -960 423588 480 423678
rect 2957 423675 3023 423678
rect 583520 416530 584960 416620
rect 583342 416470 584960 416530
rect 348918 415652 348924 415716
rect 348988 415714 348994 415716
rect 348988 415654 354690 415714
rect 348988 415652 348994 415654
rect 354630 415578 354690 415654
rect 364382 415654 374010 415714
rect 354630 415518 364258 415578
rect 364198 415442 364258 415518
rect 364382 415442 364442 415654
rect 373950 415578 374010 415654
rect 383702 415654 393330 415714
rect 373950 415518 383578 415578
rect 364198 415382 364442 415442
rect 383518 415442 383578 415518
rect 383702 415442 383762 415654
rect 393270 415578 393330 415654
rect 403022 415654 412650 415714
rect 393270 415518 402898 415578
rect 383518 415382 383762 415442
rect 402838 415442 402898 415518
rect 403022 415442 403082 415654
rect 412590 415578 412650 415654
rect 422342 415654 431970 415714
rect 412590 415518 422218 415578
rect 402838 415382 403082 415442
rect 422158 415442 422218 415518
rect 422342 415442 422402 415654
rect 431910 415578 431970 415654
rect 441662 415654 451290 415714
rect 431910 415518 441538 415578
rect 422158 415382 422402 415442
rect 441478 415442 441538 415518
rect 441662 415442 441722 415654
rect 451230 415578 451290 415654
rect 460982 415654 470610 415714
rect 451230 415518 460858 415578
rect 441478 415382 441722 415442
rect 460798 415442 460858 415518
rect 460982 415442 461042 415654
rect 470550 415578 470610 415654
rect 480302 415654 489930 415714
rect 470550 415518 480178 415578
rect 460798 415382 461042 415442
rect 480118 415442 480178 415518
rect 480302 415442 480362 415654
rect 489870 415578 489930 415654
rect 499622 415654 509250 415714
rect 489870 415518 499498 415578
rect 480118 415382 480362 415442
rect 499438 415442 499498 415518
rect 499622 415442 499682 415654
rect 509190 415578 509250 415654
rect 518942 415654 528570 415714
rect 509190 415518 518818 415578
rect 499438 415382 499682 415442
rect 518758 415442 518818 415518
rect 518942 415442 519002 415654
rect 528510 415578 528570 415654
rect 538262 415654 547890 415714
rect 528510 415518 538138 415578
rect 518758 415382 519002 415442
rect 538078 415442 538138 415518
rect 538262 415442 538322 415654
rect 547830 415578 547890 415654
rect 557582 415654 567210 415714
rect 547830 415518 557458 415578
rect 538078 415382 538322 415442
rect 557398 415442 557458 415518
rect 557582 415442 557642 415654
rect 567150 415578 567210 415654
rect 583342 415578 583402 416470
rect 583520 416380 584960 416470
rect 567150 415518 576778 415578
rect 557398 415382 557642 415442
rect 576718 415442 576778 415518
rect 576902 415518 583402 415578
rect 576902 415442 576962 415518
rect 576718 415382 576962 415442
rect -960 409172 480 409412
rect 579797 404834 579863 404837
rect 583520 404834 584960 404924
rect 579797 404832 584960 404834
rect 579797 404776 579802 404832
rect 579858 404776 584960 404832
rect 579797 404774 584960 404776
rect 579797 404771 579863 404774
rect 583520 404684 584960 404774
rect -960 395042 480 395132
rect 3049 395042 3115 395045
rect -960 395040 3115 395042
rect -960 394984 3054 395040
rect 3110 394984 3115 395040
rect -960 394982 3115 394984
rect -960 394892 480 394982
rect 3049 394979 3115 394982
rect 583520 393002 584960 393092
rect 583342 392942 584960 393002
rect 348734 392260 348740 392324
rect 348804 392322 348810 392324
rect 348804 392262 354690 392322
rect 348804 392260 348810 392262
rect 354630 392186 354690 392262
rect 364382 392262 374010 392322
rect 354630 392126 364258 392186
rect 364198 392050 364258 392126
rect 364382 392050 364442 392262
rect 373950 392186 374010 392262
rect 383702 392262 393330 392322
rect 373950 392126 383578 392186
rect 364198 391990 364442 392050
rect 383518 392050 383578 392126
rect 383702 392050 383762 392262
rect 393270 392186 393330 392262
rect 403022 392262 412650 392322
rect 393270 392126 402898 392186
rect 383518 391990 383762 392050
rect 402838 392050 402898 392126
rect 403022 392050 403082 392262
rect 412590 392186 412650 392262
rect 422342 392262 431970 392322
rect 412590 392126 422218 392186
rect 402838 391990 403082 392050
rect 422158 392050 422218 392126
rect 422342 392050 422402 392262
rect 431910 392186 431970 392262
rect 441662 392262 451290 392322
rect 431910 392126 441538 392186
rect 422158 391990 422402 392050
rect 441478 392050 441538 392126
rect 441662 392050 441722 392262
rect 451230 392186 451290 392262
rect 460982 392262 470610 392322
rect 451230 392126 460858 392186
rect 441478 391990 441722 392050
rect 460798 392050 460858 392126
rect 460982 392050 461042 392262
rect 470550 392186 470610 392262
rect 480302 392262 489930 392322
rect 470550 392126 480178 392186
rect 460798 391990 461042 392050
rect 480118 392050 480178 392126
rect 480302 392050 480362 392262
rect 489870 392186 489930 392262
rect 499622 392262 509250 392322
rect 489870 392126 499498 392186
rect 480118 391990 480362 392050
rect 499438 392050 499498 392126
rect 499622 392050 499682 392262
rect 509190 392186 509250 392262
rect 518942 392262 528570 392322
rect 509190 392126 518818 392186
rect 499438 391990 499682 392050
rect 518758 392050 518818 392126
rect 518942 392050 519002 392262
rect 528510 392186 528570 392262
rect 538262 392262 547890 392322
rect 528510 392126 538138 392186
rect 518758 391990 519002 392050
rect 538078 392050 538138 392126
rect 538262 392050 538322 392262
rect 547830 392186 547890 392262
rect 557582 392262 567210 392322
rect 547830 392126 557458 392186
rect 538078 391990 538322 392050
rect 557398 392050 557458 392126
rect 557582 392050 557642 392262
rect 567150 392186 567210 392262
rect 583342 392186 583402 392942
rect 583520 392852 584960 392942
rect 567150 392126 576778 392186
rect 557398 391990 557642 392050
rect 576718 392050 576778 392126
rect 576902 392126 583402 392186
rect 576902 392050 576962 392126
rect 576718 391990 576962 392050
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 3141 380626 3207 380629
rect -960 380624 3207 380626
rect -960 380568 3146 380624
rect 3202 380568 3207 380624
rect -960 380566 3207 380568
rect -960 380476 480 380566
rect 3141 380563 3207 380566
rect 583520 369610 584960 369700
rect 583342 369550 584960 369610
rect 348550 368732 348556 368796
rect 348620 368794 348626 368796
rect 348620 368734 354690 368794
rect 348620 368732 348626 368734
rect 354630 368658 354690 368734
rect 364382 368734 374010 368794
rect 354630 368598 364258 368658
rect 364198 368522 364258 368598
rect 364382 368522 364442 368734
rect 373950 368658 374010 368734
rect 383702 368734 393330 368794
rect 373950 368598 383578 368658
rect 364198 368462 364442 368522
rect 383518 368522 383578 368598
rect 383702 368522 383762 368734
rect 393270 368658 393330 368734
rect 403022 368734 412650 368794
rect 393270 368598 402898 368658
rect 383518 368462 383762 368522
rect 402838 368522 402898 368598
rect 403022 368522 403082 368734
rect 412590 368658 412650 368734
rect 422342 368734 431970 368794
rect 412590 368598 422218 368658
rect 402838 368462 403082 368522
rect 422158 368522 422218 368598
rect 422342 368522 422402 368734
rect 431910 368658 431970 368734
rect 441662 368734 451290 368794
rect 431910 368598 441538 368658
rect 422158 368462 422402 368522
rect 441478 368522 441538 368598
rect 441662 368522 441722 368734
rect 451230 368658 451290 368734
rect 460982 368734 470610 368794
rect 451230 368598 460858 368658
rect 441478 368462 441722 368522
rect 460798 368522 460858 368598
rect 460982 368522 461042 368734
rect 470550 368658 470610 368734
rect 480302 368734 489930 368794
rect 470550 368598 480178 368658
rect 460798 368462 461042 368522
rect 480118 368522 480178 368598
rect 480302 368522 480362 368734
rect 489870 368658 489930 368734
rect 499622 368734 509250 368794
rect 489870 368598 499498 368658
rect 480118 368462 480362 368522
rect 499438 368522 499498 368598
rect 499622 368522 499682 368734
rect 509190 368658 509250 368734
rect 518942 368734 528570 368794
rect 509190 368598 518818 368658
rect 499438 368462 499682 368522
rect 518758 368522 518818 368598
rect 518942 368522 519002 368734
rect 528510 368658 528570 368734
rect 538262 368734 547890 368794
rect 528510 368598 538138 368658
rect 518758 368462 519002 368522
rect 538078 368522 538138 368598
rect 538262 368522 538322 368734
rect 547830 368658 547890 368734
rect 557582 368734 567210 368794
rect 547830 368598 557458 368658
rect 538078 368462 538322 368522
rect 557398 368522 557458 368598
rect 557582 368522 557642 368734
rect 567150 368658 567210 368734
rect 583342 368658 583402 369550
rect 583520 369460 584960 369550
rect 567150 368598 576778 368658
rect 557398 368462 557642 368522
rect 576718 368522 576778 368598
rect 576902 368598 583402 368658
rect 576902 368522 576962 368598
rect 576718 368462 576962 368522
rect -960 366210 480 366300
rect 3233 366210 3299 366213
rect -960 366208 3299 366210
rect -960 366152 3238 366208
rect 3294 366152 3299 366208
rect -960 366150 3299 366152
rect -960 366060 480 366150
rect 3233 366147 3299 366150
rect 579889 357914 579955 357917
rect 583520 357914 584960 358004
rect 579889 357912 584960 357914
rect 579889 357856 579894 357912
rect 579950 357856 584960 357912
rect 579889 357854 584960 357856
rect 579889 357851 579955 357854
rect 583520 357764 584960 357854
rect -960 351780 480 352020
rect 583520 346082 584960 346172
rect 583342 346022 584960 346082
rect 348366 345340 348372 345404
rect 348436 345402 348442 345404
rect 348436 345342 354690 345402
rect 348436 345340 348442 345342
rect 354630 345266 354690 345342
rect 364382 345342 374010 345402
rect 354630 345206 364258 345266
rect 364198 345130 364258 345206
rect 364382 345130 364442 345342
rect 373950 345266 374010 345342
rect 383702 345342 393330 345402
rect 373950 345206 383578 345266
rect 364198 345070 364442 345130
rect 383518 345130 383578 345206
rect 383702 345130 383762 345342
rect 393270 345266 393330 345342
rect 403022 345342 412650 345402
rect 393270 345206 402898 345266
rect 383518 345070 383762 345130
rect 402838 345130 402898 345206
rect 403022 345130 403082 345342
rect 412590 345266 412650 345342
rect 422342 345342 431970 345402
rect 412590 345206 422218 345266
rect 402838 345070 403082 345130
rect 422158 345130 422218 345206
rect 422342 345130 422402 345342
rect 431910 345266 431970 345342
rect 441662 345342 451290 345402
rect 431910 345206 441538 345266
rect 422158 345070 422402 345130
rect 441478 345130 441538 345206
rect 441662 345130 441722 345342
rect 451230 345266 451290 345342
rect 460982 345342 470610 345402
rect 451230 345206 460858 345266
rect 441478 345070 441722 345130
rect 460798 345130 460858 345206
rect 460982 345130 461042 345342
rect 470550 345266 470610 345342
rect 480302 345342 489930 345402
rect 470550 345206 480178 345266
rect 460798 345070 461042 345130
rect 480118 345130 480178 345206
rect 480302 345130 480362 345342
rect 489870 345266 489930 345342
rect 499622 345342 509250 345402
rect 489870 345206 499498 345266
rect 480118 345070 480362 345130
rect 499438 345130 499498 345206
rect 499622 345130 499682 345342
rect 509190 345266 509250 345342
rect 518942 345342 528570 345402
rect 509190 345206 518818 345266
rect 499438 345070 499682 345130
rect 518758 345130 518818 345206
rect 518942 345130 519002 345342
rect 528510 345266 528570 345342
rect 538262 345342 547890 345402
rect 528510 345206 538138 345266
rect 518758 345070 519002 345130
rect 538078 345130 538138 345206
rect 538262 345130 538322 345342
rect 547830 345266 547890 345342
rect 557582 345342 567210 345402
rect 547830 345206 557458 345266
rect 538078 345070 538322 345130
rect 557398 345130 557458 345206
rect 557582 345130 557642 345342
rect 567150 345266 567210 345342
rect 583342 345266 583402 346022
rect 583520 345932 584960 346022
rect 567150 345206 576778 345266
rect 557398 345070 557642 345130
rect 576718 345130 576778 345206
rect 576902 345206 583402 345266
rect 576902 345130 576962 345206
rect 576718 345070 576962 345130
rect 266353 338194 266419 338197
rect 266353 338192 266554 338194
rect 266353 338136 266358 338192
rect 266414 338136 266554 338192
rect 266353 338134 266554 338136
rect 266353 338131 266419 338134
rect 231209 338058 231275 338061
rect 231577 338058 231643 338061
rect 266494 338060 266554 338134
rect 231209 338056 231643 338058
rect 231209 338000 231214 338056
rect 231270 338000 231582 338056
rect 231638 338000 231643 338056
rect 231209 337998 231643 338000
rect 231209 337995 231275 337998
rect 231577 337995 231643 337998
rect 266486 337996 266492 338060
rect 266556 337996 266562 338060
rect 37181 337786 37247 337789
rect 331305 337786 331371 337789
rect 37181 337784 331371 337786
rect 37181 337728 37186 337784
rect 37242 337728 331310 337784
rect 331366 337728 331371 337784
rect 37181 337726 331371 337728
rect 37181 337723 37247 337726
rect 331305 337723 331371 337726
rect 22001 337650 22067 337653
rect 328177 337650 328243 337653
rect 22001 337648 328243 337650
rect -960 337514 480 337604
rect 22001 337592 22006 337648
rect 22062 337592 328182 337648
rect 328238 337592 328243 337648
rect 22001 337590 328243 337592
rect 22001 337587 22067 337590
rect 328177 337587 328243 337590
rect 3325 337514 3391 337517
rect -960 337512 3391 337514
rect -960 337456 3330 337512
rect 3386 337456 3391 337512
rect -960 337454 3391 337456
rect -960 337364 480 337454
rect 3325 337451 3391 337454
rect 12341 337514 12407 337517
rect 326153 337514 326219 337517
rect 12341 337512 326219 337514
rect 12341 337456 12346 337512
rect 12402 337456 326158 337512
rect 326214 337456 326219 337512
rect 12341 337454 326219 337456
rect 12341 337451 12407 337454
rect 326153 337451 326219 337454
rect 10961 337378 11027 337381
rect 325969 337378 326035 337381
rect 10961 337376 326035 337378
rect 10961 337320 10966 337376
rect 11022 337320 325974 337376
rect 326030 337320 326035 337376
rect 10961 337318 326035 337320
rect 10961 337315 11027 337318
rect 325969 337315 326035 337318
rect 322013 337242 322079 337245
rect 323945 337242 324011 337245
rect 322013 337240 324011 337242
rect 322013 337184 322018 337240
rect 322074 337184 323950 337240
rect 324006 337184 324011 337240
rect 322013 337182 324011 337184
rect 322013 337179 322079 337182
rect 323945 337179 324011 337182
rect 262949 336970 263015 336973
rect 262630 336968 263015 336970
rect 262630 336912 262954 336968
rect 263010 336912 263015 336968
rect 262630 336910 263015 336912
rect 262630 336834 262690 336910
rect 262949 336907 263015 336910
rect 272241 336970 272307 336973
rect 305177 336970 305243 336973
rect 272241 336968 272580 336970
rect 272241 336912 272246 336968
rect 272302 336912 272580 336968
rect 272241 336910 272580 336912
rect 272241 336907 272307 336910
rect 272520 336837 272580 336910
rect 305177 336968 305562 336970
rect 305177 336912 305182 336968
rect 305238 336912 305562 336968
rect 305177 336910 305562 336912
rect 305177 336907 305243 336910
rect 262765 336834 262831 336837
rect 262630 336832 262831 336834
rect 262630 336776 262770 336832
rect 262826 336776 262831 336832
rect 262630 336774 262831 336776
rect 262765 336771 262831 336774
rect 272517 336832 272583 336837
rect 272517 336776 272522 336832
rect 272578 336776 272583 336832
rect 272517 336771 272583 336776
rect 305361 336834 305427 336837
rect 305502 336834 305562 336910
rect 305361 336832 305562 336834
rect 305361 336776 305366 336832
rect 305422 336776 305562 336832
rect 305361 336774 305562 336776
rect 305361 336771 305427 336774
rect 272333 336698 272399 336701
rect 272517 336698 272583 336701
rect 272333 336696 272583 336698
rect 272333 336640 272338 336696
rect 272394 336640 272522 336696
rect 272578 336640 272583 336696
rect 272333 336638 272583 336640
rect 272333 336635 272399 336638
rect 272517 336635 272583 336638
rect 318149 335338 318215 335341
rect 318425 335338 318491 335341
rect 318149 335336 318491 335338
rect 318149 335280 318154 335336
rect 318210 335280 318430 335336
rect 318486 335280 318491 335336
rect 318149 335278 318491 335280
rect 318149 335275 318215 335278
rect 318425 335275 318491 335278
rect 330753 335338 330819 335341
rect 330937 335338 331003 335341
rect 330753 335336 331003 335338
rect 330753 335280 330758 335336
rect 330814 335280 330942 335336
rect 330998 335280 331003 335336
rect 330753 335278 331003 335280
rect 330753 335275 330819 335278
rect 330937 335275 331003 335278
rect 583520 334236 584960 334476
rect 255037 328674 255103 328677
rect 254534 328672 255103 328674
rect 254534 328616 255042 328672
rect 255098 328616 255103 328672
rect 254534 328614 255103 328616
rect 254534 328538 254594 328614
rect 255037 328611 255103 328614
rect 254669 328538 254735 328541
rect 254534 328536 254735 328538
rect 254534 328480 254674 328536
rect 254730 328480 254735 328536
rect 254534 328478 254735 328480
rect 254669 328475 254735 328478
rect 256693 328538 256759 328541
rect 257061 328538 257127 328541
rect 256693 328536 257127 328538
rect 256693 328480 256698 328536
rect 256754 328480 257066 328536
rect 257122 328480 257127 328536
rect 256693 328478 257127 328480
rect 256693 328475 256759 328478
rect 257061 328475 257127 328478
rect 266486 328476 266492 328540
rect 266556 328476 266562 328540
rect 266494 328402 266554 328476
rect 266905 328402 266971 328405
rect 266494 328400 266971 328402
rect 266494 328344 266910 328400
rect 266966 328344 266971 328400
rect 266494 328342 266971 328344
rect 266905 328339 266971 328342
rect 319437 325682 319503 325685
rect 319621 325682 319687 325685
rect 319437 325680 319687 325682
rect 319437 325624 319442 325680
rect 319498 325624 319626 325680
rect 319682 325624 319687 325680
rect 319437 325622 319687 325624
rect 319437 325619 319503 325622
rect 319621 325619 319687 325622
rect -960 323098 480 323188
rect 2773 323098 2839 323101
rect -960 323096 2839 323098
rect -960 323040 2778 323096
rect 2834 323040 2839 323096
rect -960 323038 2839 323040
rect -960 322948 480 323038
rect 2773 323035 2839 323038
rect 579981 322690 580047 322693
rect 583520 322690 584960 322780
rect 579981 322688 584960 322690
rect 579981 322632 579986 322688
rect 580042 322632 584960 322688
rect 579981 322630 584960 322632
rect 579981 322627 580047 322630
rect 583520 322540 584960 322630
rect 371877 310994 371943 310997
rect 367142 310992 371943 310994
rect 367142 310936 371882 310992
rect 371938 310936 371943 310992
rect 367142 310934 371943 310936
rect 344318 310660 344324 310724
rect 344388 310722 344394 310724
rect 350441 310722 350507 310725
rect 344388 310720 350507 310722
rect 344388 310664 350446 310720
rect 350502 310664 350507 310720
rect 344388 310662 350507 310664
rect 344388 310660 344394 310662
rect 350441 310659 350507 310662
rect 367001 310722 367067 310725
rect 367142 310722 367202 310934
rect 371877 310931 371943 310934
rect 376702 310796 376708 310860
rect 376772 310858 376778 310860
rect 583520 310858 584960 310948
rect 376772 310798 393330 310858
rect 376772 310796 376778 310798
rect 367001 310720 367202 310722
rect 367001 310664 367006 310720
rect 367062 310664 367202 310720
rect 367001 310662 367202 310664
rect 393270 310722 393330 310798
rect 403022 310798 412650 310858
rect 393270 310662 402898 310722
rect 367001 310659 367067 310662
rect 350625 310586 350691 310589
rect 357382 310586 357388 310588
rect 350625 310584 357388 310586
rect 350625 310528 350630 310584
rect 350686 310528 357388 310584
rect 350625 310526 357388 310528
rect 350625 310523 350691 310526
rect 357382 310524 357388 310526
rect 357452 310524 357458 310588
rect 371877 310586 371943 310589
rect 376702 310586 376708 310588
rect 371877 310584 376708 310586
rect 371877 310528 371882 310584
rect 371938 310528 376708 310584
rect 371877 310526 376708 310528
rect 371877 310523 371943 310526
rect 376702 310524 376708 310526
rect 376772 310524 376778 310588
rect 402838 310586 402898 310662
rect 403022 310586 403082 310798
rect 412590 310722 412650 310798
rect 422342 310798 431970 310858
rect 412590 310662 422218 310722
rect 402838 310526 403082 310586
rect 422158 310586 422218 310662
rect 422342 310586 422402 310798
rect 431910 310722 431970 310798
rect 441662 310798 451290 310858
rect 431910 310662 441538 310722
rect 422158 310526 422402 310586
rect 441478 310586 441538 310662
rect 441662 310586 441722 310798
rect 451230 310722 451290 310798
rect 460982 310798 470610 310858
rect 451230 310662 460858 310722
rect 441478 310526 441722 310586
rect 460798 310586 460858 310662
rect 460982 310586 461042 310798
rect 470550 310722 470610 310798
rect 480302 310798 489930 310858
rect 470550 310662 480178 310722
rect 460798 310526 461042 310586
rect 480118 310586 480178 310662
rect 480302 310586 480362 310798
rect 489870 310722 489930 310798
rect 499622 310798 509250 310858
rect 489870 310662 499498 310722
rect 480118 310526 480362 310586
rect 499438 310586 499498 310662
rect 499622 310586 499682 310798
rect 509190 310722 509250 310798
rect 518942 310798 528570 310858
rect 509190 310662 518818 310722
rect 499438 310526 499682 310586
rect 518758 310586 518818 310662
rect 518942 310586 519002 310798
rect 528510 310722 528570 310798
rect 538262 310798 547890 310858
rect 528510 310662 538138 310722
rect 518758 310526 519002 310586
rect 538078 310586 538138 310662
rect 538262 310586 538322 310798
rect 547830 310722 547890 310798
rect 557582 310798 567210 310858
rect 547830 310662 557458 310722
rect 538078 310526 538322 310586
rect 557398 310586 557458 310662
rect 557582 310586 557642 310798
rect 567150 310722 567210 310798
rect 583342 310798 584960 310858
rect 583342 310722 583402 310798
rect 567150 310662 576778 310722
rect 557398 310526 557642 310586
rect 576718 310586 576778 310662
rect 576902 310662 583402 310722
rect 583520 310708 584960 310798
rect 576902 310586 576962 310662
rect 576718 310526 576962 310586
rect 357382 310252 357388 310316
rect 357452 310314 357458 310316
rect 367001 310314 367067 310317
rect 357452 310312 367067 310314
rect 357452 310256 367006 310312
rect 367062 310256 367067 310312
rect 357452 310254 367067 310256
rect 357452 310252 357458 310254
rect 367001 310251 367067 310254
rect -960 308818 480 308908
rect 4061 308818 4127 308821
rect -960 308816 4127 308818
rect -960 308760 4066 308816
rect 4122 308760 4127 308816
rect -960 308758 4127 308760
rect -960 308668 480 308758
rect 4061 308755 4127 308758
rect 580073 299162 580139 299165
rect 583520 299162 584960 299252
rect 580073 299160 584960 299162
rect 580073 299104 580078 299160
rect 580134 299104 584960 299160
rect 580073 299102 584960 299104
rect 580073 299099 580139 299102
rect 583520 299012 584960 299102
rect 258809 298074 258875 298077
rect 258766 298072 258875 298074
rect 258766 298016 258814 298072
rect 258870 298016 258875 298072
rect 258766 298011 258875 298016
rect 329005 298074 329071 298077
rect 329189 298074 329255 298077
rect 329005 298072 329255 298074
rect 329005 298016 329010 298072
rect 329066 298016 329194 298072
rect 329250 298016 329255 298072
rect 329005 298014 329255 298016
rect 329005 298011 329071 298014
rect 329189 298011 329255 298014
rect 258766 297941 258826 298011
rect 258717 297936 258826 297941
rect 258717 297880 258722 297936
rect 258778 297880 258826 297936
rect 258717 297878 258826 297880
rect 258717 297875 258783 297878
rect 326245 296714 326311 296717
rect 326429 296714 326495 296717
rect 326245 296712 326495 296714
rect 326245 296656 326250 296712
rect 326306 296656 326434 296712
rect 326490 296656 326495 296712
rect 326245 296654 326495 296656
rect 326245 296651 326311 296654
rect 326429 296651 326495 296654
rect -960 294402 480 294492
rect 3969 294402 4035 294405
rect -960 294400 4035 294402
rect -960 294344 3974 294400
rect 4030 294344 4035 294400
rect -960 294342 4035 294344
rect -960 294252 480 294342
rect 3969 294339 4035 294342
rect 293125 288418 293191 288421
rect 293309 288418 293375 288421
rect 293125 288416 293375 288418
rect 293125 288360 293130 288416
rect 293186 288360 293314 288416
rect 293370 288360 293375 288416
rect 293125 288358 293375 288360
rect 293125 288355 293191 288358
rect 293309 288355 293375 288358
rect 329005 288418 329071 288421
rect 329189 288418 329255 288421
rect 329005 288416 329255 288418
rect 329005 288360 329010 288416
rect 329066 288360 329194 288416
rect 329250 288360 329255 288416
rect 329005 288358 329255 288360
rect 329005 288355 329071 288358
rect 329189 288355 329255 288358
rect 335813 288418 335879 288421
rect 335997 288418 336063 288421
rect 335813 288416 336063 288418
rect 335813 288360 335818 288416
rect 335874 288360 336002 288416
rect 336058 288360 336063 288416
rect 335813 288358 336063 288360
rect 335813 288355 335879 288358
rect 335997 288355 336063 288358
rect 583520 287316 584960 287556
rect -960 280122 480 280212
rect 2773 280122 2839 280125
rect -960 280120 2839 280122
rect -960 280064 2778 280120
rect 2834 280064 2839 280120
rect -960 280062 2839 280064
rect -960 279972 480 280062
rect 2773 280059 2839 280062
rect 107469 278762 107535 278765
rect 107653 278762 107719 278765
rect 107469 278760 107719 278762
rect 107469 278704 107474 278760
rect 107530 278704 107658 278760
rect 107714 278704 107719 278760
rect 107469 278702 107719 278704
rect 107469 278699 107535 278702
rect 107653 278699 107719 278702
rect 231945 278762 232011 278765
rect 232129 278762 232195 278765
rect 231945 278760 232195 278762
rect 231945 278704 231950 278760
rect 232006 278704 232134 278760
rect 232190 278704 232195 278760
rect 231945 278702 232195 278704
rect 231945 278699 232011 278702
rect 232129 278699 232195 278702
rect 261385 278762 261451 278765
rect 261569 278762 261635 278765
rect 261385 278760 261635 278762
rect 261385 278704 261390 278760
rect 261446 278704 261574 278760
rect 261630 278704 261635 278760
rect 261385 278702 261635 278704
rect 261385 278699 261451 278702
rect 261569 278699 261635 278702
rect 320909 278762 320975 278765
rect 321093 278762 321159 278765
rect 320909 278760 321159 278762
rect 320909 278704 320914 278760
rect 320970 278704 321098 278760
rect 321154 278704 321159 278760
rect 320909 278702 321159 278704
rect 320909 278699 320975 278702
rect 321093 278699 321159 278702
rect 319437 277402 319503 277405
rect 319621 277402 319687 277405
rect 319437 277400 319687 277402
rect 319437 277344 319442 277400
rect 319498 277344 319626 277400
rect 319682 277344 319687 277400
rect 319437 277342 319687 277344
rect 319437 277339 319503 277342
rect 319621 277339 319687 277342
rect 326245 277402 326311 277405
rect 326521 277402 326587 277405
rect 326245 277400 326587 277402
rect 326245 277344 326250 277400
rect 326306 277344 326526 277400
rect 326582 277344 326587 277400
rect 326245 277342 326587 277344
rect 326245 277339 326311 277342
rect 326521 277339 326587 277342
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect 340045 270738 340111 270741
rect 339910 270736 340111 270738
rect 339910 270680 340050 270736
rect 340106 270680 340111 270736
rect 339910 270678 340111 270680
rect 339910 270466 339970 270678
rect 340045 270675 340111 270678
rect 340321 270466 340387 270469
rect 339910 270464 340387 270466
rect 339910 270408 340326 270464
rect 340382 270408 340387 270464
rect 339910 270406 340387 270408
rect 340321 270403 340387 270406
rect 253013 269106 253079 269109
rect 264329 269106 264395 269109
rect 264513 269106 264579 269109
rect 253013 269104 253122 269106
rect 253013 269048 253018 269104
rect 253074 269048 253122 269104
rect 253013 269043 253122 269048
rect 264329 269104 264579 269106
rect 264329 269048 264334 269104
rect 264390 269048 264518 269104
rect 264574 269048 264579 269104
rect 264329 269046 264579 269048
rect 264329 269043 264395 269046
rect 264513 269043 264579 269046
rect 265617 269106 265683 269109
rect 265801 269106 265867 269109
rect 265617 269104 265867 269106
rect 265617 269048 265622 269104
rect 265678 269048 265806 269104
rect 265862 269048 265867 269104
rect 265617 269046 265867 269048
rect 265617 269043 265683 269046
rect 265801 269043 265867 269046
rect 293125 269106 293191 269109
rect 293309 269106 293375 269109
rect 293125 269104 293375 269106
rect 293125 269048 293130 269104
rect 293186 269048 293314 269104
rect 293370 269048 293375 269104
rect 293125 269046 293375 269048
rect 293125 269043 293191 269046
rect 293309 269043 293375 269046
rect 320909 269106 320975 269109
rect 321093 269106 321159 269109
rect 320909 269104 321159 269106
rect 320909 269048 320914 269104
rect 320970 269048 321098 269104
rect 321154 269048 321159 269104
rect 320909 269046 321159 269048
rect 320909 269043 320975 269046
rect 321093 269043 321159 269046
rect 253062 268973 253122 269043
rect 253062 268968 253171 268973
rect 253062 268912 253110 268968
rect 253166 268912 253171 268968
rect 253062 268910 253171 268912
rect 253105 268907 253171 268910
rect 246481 267882 246547 267885
rect 246757 267882 246823 267885
rect 246481 267880 246823 267882
rect 246481 267824 246486 267880
rect 246542 267824 246762 267880
rect 246818 267824 246823 267880
rect 246481 267822 246823 267824
rect 246481 267819 246547 267822
rect 246757 267819 246823 267822
rect 246297 267746 246363 267749
rect 246481 267746 246547 267749
rect 246297 267744 246547 267746
rect 246297 267688 246302 267744
rect 246358 267688 246486 267744
rect 246542 267688 246547 267744
rect 246297 267686 246547 267688
rect 246297 267683 246363 267686
rect 246481 267683 246547 267686
rect -960 265706 480 265796
rect 2773 265706 2839 265709
rect -960 265704 2839 265706
rect -960 265648 2778 265704
rect 2834 265648 2839 265704
rect -960 265646 2839 265648
rect -960 265556 480 265646
rect 2773 265643 2839 265646
rect 371877 264074 371943 264077
rect 367142 264072 371943 264074
rect 367142 264016 371882 264072
rect 371938 264016 371943 264072
rect 367142 264014 371943 264016
rect 344134 263740 344140 263804
rect 344204 263802 344210 263804
rect 350441 263802 350507 263805
rect 344204 263800 350507 263802
rect 344204 263744 350446 263800
rect 350502 263744 350507 263800
rect 344204 263742 350507 263744
rect 344204 263740 344210 263742
rect 350441 263739 350507 263742
rect 367001 263802 367067 263805
rect 367142 263802 367202 264014
rect 371877 264011 371943 264014
rect 376702 263876 376708 263940
rect 376772 263938 376778 263940
rect 583520 263938 584960 264028
rect 376772 263878 393330 263938
rect 376772 263876 376778 263878
rect 367001 263800 367202 263802
rect 367001 263744 367006 263800
rect 367062 263744 367202 263800
rect 367001 263742 367202 263744
rect 393270 263802 393330 263878
rect 403022 263878 412650 263938
rect 393270 263742 402898 263802
rect 367001 263739 367067 263742
rect 350625 263666 350691 263669
rect 357382 263666 357388 263668
rect 350625 263664 357388 263666
rect 350625 263608 350630 263664
rect 350686 263608 357388 263664
rect 350625 263606 357388 263608
rect 350625 263603 350691 263606
rect 357382 263604 357388 263606
rect 357452 263604 357458 263668
rect 371877 263666 371943 263669
rect 376702 263666 376708 263668
rect 371877 263664 376708 263666
rect 371877 263608 371882 263664
rect 371938 263608 376708 263664
rect 371877 263606 376708 263608
rect 371877 263603 371943 263606
rect 376702 263604 376708 263606
rect 376772 263604 376778 263668
rect 402838 263666 402898 263742
rect 403022 263666 403082 263878
rect 412590 263802 412650 263878
rect 422342 263878 431970 263938
rect 412590 263742 422218 263802
rect 402838 263606 403082 263666
rect 422158 263666 422218 263742
rect 422342 263666 422402 263878
rect 431910 263802 431970 263878
rect 441662 263878 451290 263938
rect 431910 263742 441538 263802
rect 422158 263606 422402 263666
rect 441478 263666 441538 263742
rect 441662 263666 441722 263878
rect 451230 263802 451290 263878
rect 460982 263878 470610 263938
rect 451230 263742 460858 263802
rect 441478 263606 441722 263666
rect 460798 263666 460858 263742
rect 460982 263666 461042 263878
rect 470550 263802 470610 263878
rect 480302 263878 489930 263938
rect 470550 263742 480178 263802
rect 460798 263606 461042 263666
rect 480118 263666 480178 263742
rect 480302 263666 480362 263878
rect 489870 263802 489930 263878
rect 499622 263878 509250 263938
rect 489870 263742 499498 263802
rect 480118 263606 480362 263666
rect 499438 263666 499498 263742
rect 499622 263666 499682 263878
rect 509190 263802 509250 263878
rect 518942 263878 528570 263938
rect 509190 263742 518818 263802
rect 499438 263606 499682 263666
rect 518758 263666 518818 263742
rect 518942 263666 519002 263878
rect 528510 263802 528570 263878
rect 538262 263878 547890 263938
rect 528510 263742 538138 263802
rect 518758 263606 519002 263666
rect 538078 263666 538138 263742
rect 538262 263666 538322 263878
rect 547830 263802 547890 263878
rect 557582 263878 567210 263938
rect 547830 263742 557458 263802
rect 538078 263606 538322 263666
rect 557398 263666 557458 263742
rect 557582 263666 557642 263878
rect 567150 263802 567210 263878
rect 583342 263878 584960 263938
rect 583342 263802 583402 263878
rect 567150 263742 576778 263802
rect 557398 263606 557642 263666
rect 576718 263666 576778 263742
rect 576902 263742 583402 263802
rect 583520 263788 584960 263878
rect 576902 263666 576962 263742
rect 576718 263606 576962 263666
rect 357382 263332 357388 263396
rect 357452 263394 357458 263396
rect 367001 263394 367067 263397
rect 357452 263392 367067 263394
rect 357452 263336 367006 263392
rect 367062 263336 367067 263392
rect 357452 263334 367067 263336
rect 357452 263332 357458 263334
rect 367001 263331 367067 263334
rect 107469 259450 107535 259453
rect 107653 259450 107719 259453
rect 107469 259448 107719 259450
rect 107469 259392 107474 259448
rect 107530 259392 107658 259448
rect 107714 259392 107719 259448
rect 107469 259390 107719 259392
rect 107469 259387 107535 259390
rect 107653 259387 107719 259390
rect 320909 259450 320975 259453
rect 321093 259450 321159 259453
rect 322289 259450 322355 259453
rect 320909 259448 321159 259450
rect 320909 259392 320914 259448
rect 320970 259392 321098 259448
rect 321154 259392 321159 259448
rect 320909 259390 321159 259392
rect 320909 259387 320975 259390
rect 321093 259387 321159 259390
rect 322246 259448 322355 259450
rect 322246 259392 322294 259448
rect 322350 259392 322355 259448
rect 322246 259387 322355 259392
rect 345381 259450 345447 259453
rect 345565 259450 345631 259453
rect 345381 259448 345631 259450
rect 345381 259392 345386 259448
rect 345442 259392 345570 259448
rect 345626 259392 345631 259448
rect 345381 259390 345631 259392
rect 345381 259387 345447 259390
rect 345565 259387 345631 259390
rect 322246 259317 322306 259387
rect 322197 259312 322306 259317
rect 322197 259256 322202 259312
rect 322258 259256 322306 259312
rect 322197 259254 322306 259256
rect 322197 259251 322263 259254
rect 231761 258090 231827 258093
rect 231945 258090 232011 258093
rect 231761 258088 232011 258090
rect 231761 258032 231766 258088
rect 231822 258032 231950 258088
rect 232006 258032 232011 258088
rect 231761 258030 232011 258032
rect 231761 258027 231827 258030
rect 231945 258027 232011 258030
rect 244365 258090 244431 258093
rect 244641 258090 244707 258093
rect 244365 258088 244707 258090
rect 244365 258032 244370 258088
rect 244426 258032 244646 258088
rect 244702 258032 244707 258088
rect 244365 258030 244707 258032
rect 244365 258027 244431 258030
rect 244641 258027 244707 258030
rect 331581 256730 331647 256733
rect 331765 256730 331831 256733
rect 331581 256728 331831 256730
rect 331581 256672 331586 256728
rect 331642 256672 331770 256728
rect 331826 256672 331831 256728
rect 331581 256670 331831 256672
rect 331581 256667 331647 256670
rect 331765 256667 331831 256670
rect 580901 252242 580967 252245
rect 583520 252242 584960 252332
rect 580901 252240 584960 252242
rect 580901 252184 580906 252240
rect 580962 252184 584960 252240
rect 580901 252182 584960 252184
rect 580901 252179 580967 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3877 251290 3943 251293
rect -960 251288 3943 251290
rect -960 251232 3882 251288
rect 3938 251232 3943 251288
rect -960 251230 3943 251232
rect -960 251140 480 251230
rect 3877 251227 3943 251230
rect 264329 249794 264395 249797
rect 264513 249794 264579 249797
rect 264329 249792 264579 249794
rect 264329 249736 264334 249792
rect 264390 249736 264518 249792
rect 264574 249736 264579 249792
rect 264329 249734 264579 249736
rect 264329 249731 264395 249734
rect 264513 249731 264579 249734
rect 293125 249794 293191 249797
rect 293309 249794 293375 249797
rect 293125 249792 293375 249794
rect 293125 249736 293130 249792
rect 293186 249736 293314 249792
rect 293370 249736 293375 249792
rect 293125 249734 293375 249736
rect 293125 249731 293191 249734
rect 293309 249731 293375 249734
rect 320909 249794 320975 249797
rect 321093 249794 321159 249797
rect 320909 249792 321159 249794
rect 320909 249736 320914 249792
rect 320970 249736 321098 249792
rect 321154 249736 321159 249792
rect 320909 249734 321159 249736
rect 320909 249731 320975 249734
rect 321093 249731 321159 249734
rect 260189 248434 260255 248437
rect 260373 248434 260439 248437
rect 260189 248432 260439 248434
rect 260189 248376 260194 248432
rect 260250 248376 260378 248432
rect 260434 248376 260439 248432
rect 260189 248374 260439 248376
rect 260189 248371 260255 248374
rect 260373 248371 260439 248374
rect 265617 248434 265683 248437
rect 265801 248434 265867 248437
rect 265617 248432 265867 248434
rect 265617 248376 265622 248432
rect 265678 248376 265806 248432
rect 265862 248376 265867 248432
rect 265617 248374 265867 248376
rect 265617 248371 265683 248374
rect 265801 248371 265867 248374
rect 322105 248434 322171 248437
rect 322289 248434 322355 248437
rect 322105 248432 322355 248434
rect 322105 248376 322110 248432
rect 322166 248376 322294 248432
rect 322350 248376 322355 248432
rect 322105 248374 322355 248376
rect 322105 248371 322171 248374
rect 322289 248371 322355 248374
rect 330569 247346 330635 247349
rect 330526 247344 330635 247346
rect 330526 247288 330574 247344
rect 330630 247288 330635 247344
rect 330526 247283 330635 247288
rect 330526 247077 330586 247283
rect 333237 247210 333303 247213
rect 333237 247208 333346 247210
rect 333237 247152 333242 247208
rect 333298 247152 333346 247208
rect 333237 247147 333346 247152
rect 333286 247077 333346 247147
rect 330526 247072 330635 247077
rect 330526 247016 330574 247072
rect 330630 247016 330635 247072
rect 330526 247014 330635 247016
rect 330569 247011 330635 247014
rect 333237 247072 333346 247077
rect 333237 247016 333242 247072
rect 333298 247016 333346 247072
rect 333237 247014 333346 247016
rect 333237 247011 333303 247014
rect 107469 241770 107535 241773
rect 107334 241768 107535 241770
rect 107334 241712 107474 241768
rect 107530 241712 107535 241768
rect 107334 241710 107535 241712
rect 107334 241634 107394 241710
rect 107469 241707 107535 241710
rect 107469 241634 107535 241637
rect 107334 241632 107535 241634
rect 107334 241576 107474 241632
rect 107530 241576 107535 241632
rect 107334 241574 107535 241576
rect 107469 241571 107535 241574
rect 231209 241498 231275 241501
rect 231393 241498 231459 241501
rect 231209 241496 231459 241498
rect 231209 241440 231214 241496
rect 231270 241440 231398 241496
rect 231454 241440 231459 241496
rect 231209 241438 231459 241440
rect 231209 241435 231275 241438
rect 231393 241435 231459 241438
rect 583520 240396 584960 240636
rect 107469 240138 107535 240141
rect 107653 240138 107719 240141
rect 107469 240136 107719 240138
rect 107469 240080 107474 240136
rect 107530 240080 107658 240136
rect 107714 240080 107719 240136
rect 107469 240078 107719 240080
rect 107469 240075 107535 240078
rect 107653 240075 107719 240078
rect 232313 240138 232379 240141
rect 232589 240138 232655 240141
rect 232313 240136 232655 240138
rect 232313 240080 232318 240136
rect 232374 240080 232594 240136
rect 232650 240080 232655 240136
rect 232313 240078 232655 240080
rect 232313 240075 232379 240078
rect 232589 240075 232655 240078
rect 237833 240138 237899 240141
rect 238017 240138 238083 240141
rect 237833 240136 238083 240138
rect 237833 240080 237838 240136
rect 237894 240080 238022 240136
rect 238078 240080 238083 240136
rect 237833 240078 238083 240080
rect 237833 240075 237899 240078
rect 238017 240075 238083 240078
rect 240501 240138 240567 240141
rect 240685 240138 240751 240141
rect 240501 240136 240751 240138
rect 240501 240080 240506 240136
rect 240562 240080 240690 240136
rect 240746 240080 240751 240136
rect 240501 240078 240751 240080
rect 240501 240075 240567 240078
rect 240685 240075 240751 240078
rect 244181 240138 244247 240141
rect 244365 240138 244431 240141
rect 244181 240136 244431 240138
rect 244181 240080 244186 240136
rect 244242 240080 244370 240136
rect 244426 240080 244431 240136
rect 244181 240078 244431 240080
rect 244181 240075 244247 240078
rect 244365 240075 244431 240078
rect 320909 240138 320975 240141
rect 321093 240138 321159 240141
rect 320909 240136 321159 240138
rect 320909 240080 320914 240136
rect 320970 240080 321098 240136
rect 321154 240080 321159 240136
rect 320909 240078 321159 240080
rect 320909 240075 320975 240078
rect 321093 240075 321159 240078
rect 335813 238778 335879 238781
rect 335997 238778 336063 238781
rect 335813 238776 336063 238778
rect 335813 238720 335818 238776
rect 335874 238720 336002 238776
rect 336058 238720 336063 238776
rect 335813 238718 336063 238720
rect 335813 238715 335879 238718
rect 335997 238715 336063 238718
rect 331765 237418 331831 237421
rect 331949 237418 332015 237421
rect 331765 237416 332015 237418
rect 331765 237360 331770 237416
rect 331826 237360 331954 237416
rect 332010 237360 332015 237416
rect 331765 237358 332015 237360
rect 331765 237355 331831 237358
rect 331949 237355 332015 237358
rect 333237 237418 333303 237421
rect 333421 237418 333487 237421
rect 333237 237416 333487 237418
rect 333237 237360 333242 237416
rect 333298 237360 333426 237416
rect 333482 237360 333487 237416
rect 333237 237358 333487 237360
rect 333237 237355 333303 237358
rect 333421 237355 333487 237358
rect -960 237010 480 237100
rect 2773 237010 2839 237013
rect -960 237008 2839 237010
rect -960 236952 2778 237008
rect 2834 236952 2839 237008
rect -960 236950 2839 236952
rect -960 236860 480 236950
rect 2773 236947 2839 236950
rect 100661 231842 100727 231845
rect 100845 231842 100911 231845
rect 100661 231840 100911 231842
rect 100661 231784 100666 231840
rect 100722 231784 100850 231840
rect 100906 231784 100911 231840
rect 100661 231782 100911 231784
rect 100661 231779 100727 231782
rect 100845 231779 100911 231782
rect 258625 230618 258691 230621
rect 258625 230616 258826 230618
rect 258625 230560 258630 230616
rect 258686 230560 258826 230616
rect 258625 230558 258826 230560
rect 258625 230555 258691 230558
rect 258766 230485 258826 230558
rect 253013 230482 253079 230485
rect 253289 230482 253355 230485
rect 253013 230480 253355 230482
rect 253013 230424 253018 230480
rect 253074 230424 253294 230480
rect 253350 230424 253355 230480
rect 253013 230422 253355 230424
rect 253013 230419 253079 230422
rect 253289 230419 253355 230422
rect 258717 230480 258826 230485
rect 258717 230424 258722 230480
rect 258778 230424 258826 230480
rect 258717 230422 258826 230424
rect 293125 230482 293191 230485
rect 293309 230482 293375 230485
rect 293125 230480 293375 230482
rect 293125 230424 293130 230480
rect 293186 230424 293314 230480
rect 293370 230424 293375 230480
rect 293125 230422 293375 230424
rect 258717 230419 258783 230422
rect 293125 230419 293191 230422
rect 293309 230419 293375 230422
rect 320909 230482 320975 230485
rect 321093 230482 321159 230485
rect 320909 230480 321159 230482
rect 320909 230424 320914 230480
rect 320970 230424 321098 230480
rect 321154 230424 321159 230480
rect 320909 230422 321159 230424
rect 320909 230419 320975 230422
rect 321093 230419 321159 230422
rect 339953 230482 340019 230485
rect 340137 230482 340203 230485
rect 339953 230480 340203 230482
rect 339953 230424 339958 230480
rect 340014 230424 340142 230480
rect 340198 230424 340203 230480
rect 339953 230422 340203 230424
rect 339953 230419 340019 230422
rect 340137 230419 340203 230422
rect 265617 229122 265683 229125
rect 265801 229122 265867 229125
rect 265617 229120 265867 229122
rect 265617 229064 265622 229120
rect 265678 229064 265806 229120
rect 265862 229064 265867 229120
rect 265617 229062 265867 229064
rect 265617 229059 265683 229062
rect 265801 229059 265867 229062
rect 319437 229122 319503 229125
rect 319621 229122 319687 229125
rect 319437 229120 319687 229122
rect 319437 229064 319442 229120
rect 319498 229064 319626 229120
rect 319682 229064 319687 229120
rect 319437 229062 319687 229064
rect 319437 229059 319503 229062
rect 319621 229059 319687 229062
rect 322105 229122 322171 229125
rect 322289 229122 322355 229125
rect 322105 229120 322355 229122
rect 322105 229064 322110 229120
rect 322166 229064 322294 229120
rect 322350 229064 322355 229120
rect 322105 229062 322355 229064
rect 322105 229059 322171 229062
rect 322289 229059 322355 229062
rect 580809 228850 580875 228853
rect 583520 228850 584960 228940
rect 580809 228848 584960 228850
rect 580809 228792 580814 228848
rect 580870 228792 584960 228848
rect 580809 228790 584960 228792
rect 580809 228787 580875 228790
rect 583520 228700 584960 228790
rect -960 222594 480 222684
rect 2773 222594 2839 222597
rect -960 222592 2839 222594
rect -960 222536 2778 222592
rect 2834 222536 2839 222592
rect -960 222534 2839 222536
rect -960 222444 480 222534
rect 2773 222531 2839 222534
rect 231209 222186 231275 222189
rect 231393 222186 231459 222189
rect 231209 222184 231459 222186
rect 231209 222128 231214 222184
rect 231270 222128 231398 222184
rect 231454 222128 231459 222184
rect 231209 222126 231459 222128
rect 231209 222123 231275 222126
rect 231393 222123 231459 222126
rect 107469 220826 107535 220829
rect 107653 220826 107719 220829
rect 107469 220824 107719 220826
rect 107469 220768 107474 220824
rect 107530 220768 107658 220824
rect 107714 220768 107719 220824
rect 107469 220766 107719 220768
rect 107469 220763 107535 220766
rect 107653 220763 107719 220766
rect 232037 220828 232103 220829
rect 232037 220824 232084 220828
rect 232148 220826 232154 220828
rect 232313 220826 232379 220829
rect 232773 220826 232839 220829
rect 232037 220768 232042 220824
rect 232037 220764 232084 220768
rect 232148 220766 232194 220826
rect 232313 220824 232839 220826
rect 232313 220768 232318 220824
rect 232374 220768 232778 220824
rect 232834 220768 232839 220824
rect 232313 220766 232839 220768
rect 232148 220764 232154 220766
rect 232037 220763 232103 220764
rect 232313 220763 232379 220766
rect 232773 220763 232839 220766
rect 240501 220826 240567 220829
rect 240685 220826 240751 220829
rect 240501 220824 240751 220826
rect 240501 220768 240506 220824
rect 240562 220768 240690 220824
rect 240746 220768 240751 220824
rect 240501 220766 240751 220768
rect 240501 220763 240567 220766
rect 240685 220763 240751 220766
rect 293125 220826 293191 220829
rect 293309 220826 293375 220829
rect 293125 220824 293375 220826
rect 293125 220768 293130 220824
rect 293186 220768 293314 220824
rect 293370 220768 293375 220824
rect 293125 220766 293375 220768
rect 293125 220763 293191 220766
rect 293309 220763 293375 220766
rect 322105 219466 322171 219469
rect 322289 219466 322355 219469
rect 322105 219464 322355 219466
rect 322105 219408 322110 219464
rect 322166 219408 322294 219464
rect 322350 219408 322355 219464
rect 322105 219406 322355 219408
rect 322105 219403 322171 219406
rect 322289 219403 322355 219406
rect 301589 218106 301655 218109
rect 301773 218106 301839 218109
rect 301589 218104 301839 218106
rect 301589 218048 301594 218104
rect 301650 218048 301778 218104
rect 301834 218048 301839 218104
rect 301589 218046 301839 218048
rect 301589 218043 301655 218046
rect 301773 218043 301839 218046
rect 371877 217154 371943 217157
rect 367142 217152 371943 217154
rect 367142 217096 371882 217152
rect 371938 217096 371943 217152
rect 367142 217094 371943 217096
rect 342478 216820 342484 216884
rect 342548 216882 342554 216884
rect 350441 216882 350507 216885
rect 342548 216880 350507 216882
rect 342548 216824 350446 216880
rect 350502 216824 350507 216880
rect 342548 216822 350507 216824
rect 342548 216820 342554 216822
rect 350441 216819 350507 216822
rect 367001 216882 367067 216885
rect 367142 216882 367202 217094
rect 371877 217091 371943 217094
rect 376702 216956 376708 217020
rect 376772 217018 376778 217020
rect 583520 217018 584960 217108
rect 376772 216958 393330 217018
rect 376772 216956 376778 216958
rect 367001 216880 367202 216882
rect 367001 216824 367006 216880
rect 367062 216824 367202 216880
rect 367001 216822 367202 216824
rect 393270 216882 393330 216958
rect 403022 216958 412650 217018
rect 393270 216822 402898 216882
rect 367001 216819 367067 216822
rect 350625 216746 350691 216749
rect 357382 216746 357388 216748
rect 350625 216744 357388 216746
rect 350625 216688 350630 216744
rect 350686 216688 357388 216744
rect 350625 216686 357388 216688
rect 350625 216683 350691 216686
rect 357382 216684 357388 216686
rect 357452 216684 357458 216748
rect 371877 216746 371943 216749
rect 376702 216746 376708 216748
rect 371877 216744 376708 216746
rect 371877 216688 371882 216744
rect 371938 216688 376708 216744
rect 371877 216686 376708 216688
rect 371877 216683 371943 216686
rect 376702 216684 376708 216686
rect 376772 216684 376778 216748
rect 402838 216746 402898 216822
rect 403022 216746 403082 216958
rect 412590 216882 412650 216958
rect 422342 216958 431970 217018
rect 412590 216822 422218 216882
rect 402838 216686 403082 216746
rect 422158 216746 422218 216822
rect 422342 216746 422402 216958
rect 431910 216882 431970 216958
rect 441662 216958 451290 217018
rect 431910 216822 441538 216882
rect 422158 216686 422402 216746
rect 441478 216746 441538 216822
rect 441662 216746 441722 216958
rect 451230 216882 451290 216958
rect 460982 216958 470610 217018
rect 451230 216822 460858 216882
rect 441478 216686 441722 216746
rect 460798 216746 460858 216822
rect 460982 216746 461042 216958
rect 470550 216882 470610 216958
rect 480302 216958 489930 217018
rect 470550 216822 480178 216882
rect 460798 216686 461042 216746
rect 480118 216746 480178 216822
rect 480302 216746 480362 216958
rect 489870 216882 489930 216958
rect 499622 216958 509250 217018
rect 489870 216822 499498 216882
rect 480118 216686 480362 216746
rect 499438 216746 499498 216822
rect 499622 216746 499682 216958
rect 509190 216882 509250 216958
rect 518942 216958 528570 217018
rect 509190 216822 518818 216882
rect 499438 216686 499682 216746
rect 518758 216746 518818 216822
rect 518942 216746 519002 216958
rect 528510 216882 528570 216958
rect 538262 216958 547890 217018
rect 528510 216822 538138 216882
rect 518758 216686 519002 216746
rect 538078 216746 538138 216822
rect 538262 216746 538322 216958
rect 547830 216882 547890 216958
rect 557582 216958 567210 217018
rect 547830 216822 557458 216882
rect 538078 216686 538322 216746
rect 557398 216746 557458 216822
rect 557582 216746 557642 216958
rect 567150 216882 567210 216958
rect 583342 216958 584960 217018
rect 583342 216882 583402 216958
rect 567150 216822 576778 216882
rect 557398 216686 557642 216746
rect 576718 216746 576778 216822
rect 576902 216822 583402 216882
rect 583520 216868 584960 216958
rect 576902 216746 576962 216822
rect 576718 216686 576962 216746
rect 357382 216412 357388 216476
rect 357452 216474 357458 216476
rect 367001 216474 367067 216477
rect 357452 216472 367067 216474
rect 357452 216416 367006 216472
rect 367062 216416 367067 216472
rect 357452 216414 367067 216416
rect 357452 216412 357458 216414
rect 367001 216411 367067 216414
rect 330753 215386 330819 215389
rect 330937 215386 331003 215389
rect 330753 215384 331003 215386
rect 330753 215328 330758 215384
rect 330814 215328 330942 215384
rect 330998 215328 331003 215384
rect 330753 215326 331003 215328
rect 330753 215323 330819 215326
rect 330937 215323 331003 215326
rect 100661 212530 100727 212533
rect 100845 212530 100911 212533
rect 100661 212528 100911 212530
rect 100661 212472 100666 212528
rect 100722 212472 100850 212528
rect 100906 212472 100911 212528
rect 100661 212470 100911 212472
rect 100661 212467 100727 212470
rect 100845 212467 100911 212470
rect 294781 211306 294847 211309
rect 296069 211306 296135 211309
rect 294781 211304 294890 211306
rect 294781 211248 294786 211304
rect 294842 211248 294890 211304
rect 294781 211243 294890 211248
rect 296069 211304 296178 211306
rect 296069 211248 296074 211304
rect 296130 211248 296178 211304
rect 296069 211243 296178 211248
rect 294830 211173 294890 211243
rect 296118 211173 296178 211243
rect 107469 211170 107535 211173
rect 107653 211170 107719 211173
rect 232037 211172 232103 211173
rect 232037 211170 232084 211172
rect 107469 211168 107719 211170
rect 107469 211112 107474 211168
rect 107530 211112 107658 211168
rect 107714 211112 107719 211168
rect 107469 211110 107719 211112
rect 231992 211168 232084 211170
rect 231992 211112 232042 211168
rect 231992 211110 232084 211112
rect 107469 211107 107535 211110
rect 107653 211107 107719 211110
rect 232037 211108 232084 211110
rect 232148 211108 232154 211172
rect 240501 211170 240567 211173
rect 240685 211170 240751 211173
rect 240501 211168 240751 211170
rect 240501 211112 240506 211168
rect 240562 211112 240690 211168
rect 240746 211112 240751 211168
rect 240501 211110 240751 211112
rect 232037 211107 232103 211108
rect 240501 211107 240567 211110
rect 240685 211107 240751 211110
rect 253013 211170 253079 211173
rect 253197 211170 253263 211173
rect 253013 211168 253263 211170
rect 253013 211112 253018 211168
rect 253074 211112 253202 211168
rect 253258 211112 253263 211168
rect 253013 211110 253263 211112
rect 253013 211107 253079 211110
rect 253197 211107 253263 211110
rect 293125 211170 293191 211173
rect 293309 211170 293375 211173
rect 293125 211168 293375 211170
rect 293125 211112 293130 211168
rect 293186 211112 293314 211168
rect 293370 211112 293375 211168
rect 293125 211110 293375 211112
rect 293125 211107 293191 211110
rect 293309 211107 293375 211110
rect 294781 211168 294890 211173
rect 294781 211112 294786 211168
rect 294842 211112 294890 211168
rect 294781 211110 294890 211112
rect 296069 211168 296178 211173
rect 296069 211112 296074 211168
rect 296130 211112 296178 211168
rect 296069 211110 296178 211112
rect 341701 211170 341767 211173
rect 341885 211170 341951 211173
rect 341701 211168 341951 211170
rect 341701 211112 341706 211168
rect 341762 211112 341890 211168
rect 341946 211112 341951 211168
rect 341701 211110 341951 211112
rect 294781 211107 294847 211110
rect 296069 211107 296135 211110
rect 341701 211107 341767 211110
rect 341885 211107 341951 211110
rect 265617 209810 265683 209813
rect 265801 209810 265867 209813
rect 265617 209808 265867 209810
rect 265617 209752 265622 209808
rect 265678 209752 265806 209808
rect 265862 209752 265867 209808
rect 265617 209750 265867 209752
rect 265617 209747 265683 209750
rect 265801 209747 265867 209750
rect -960 208178 480 208268
rect 3785 208178 3851 208181
rect -960 208176 3851 208178
rect -960 208120 3790 208176
rect 3846 208120 3851 208176
rect -960 208118 3851 208120
rect -960 208028 480 208118
rect 3785 208115 3851 208118
rect 330753 205730 330819 205733
rect 330937 205730 331003 205733
rect 330753 205728 331003 205730
rect 330753 205672 330758 205728
rect 330814 205672 330942 205728
rect 330998 205672 331003 205728
rect 330753 205670 331003 205672
rect 330753 205667 330819 205670
rect 330937 205667 331003 205670
rect 580717 205322 580783 205325
rect 583520 205322 584960 205412
rect 580717 205320 584960 205322
rect 580717 205264 580722 205320
rect 580778 205264 584960 205320
rect 580717 205262 584960 205264
rect 580717 205259 580783 205262
rect 583520 205172 584960 205262
rect 231209 202874 231275 202877
rect 231393 202874 231459 202877
rect 231209 202872 231459 202874
rect 231209 202816 231214 202872
rect 231270 202816 231398 202872
rect 231454 202816 231459 202872
rect 231209 202814 231459 202816
rect 231209 202811 231275 202814
rect 231393 202811 231459 202814
rect 232037 202874 232103 202877
rect 232037 202872 232146 202874
rect 232037 202816 232042 202872
rect 232098 202816 232146 202872
rect 232037 202811 232146 202816
rect 232086 202741 232146 202811
rect 232086 202736 232195 202741
rect 232086 202680 232134 202736
rect 232190 202680 232195 202736
rect 232086 202678 232195 202680
rect 232129 202675 232195 202678
rect 321093 201650 321159 201653
rect 320958 201648 321159 201650
rect 320958 201592 321098 201648
rect 321154 201592 321159 201648
rect 320958 201590 321159 201592
rect 240685 201514 240751 201517
rect 240869 201514 240935 201517
rect 240685 201512 240935 201514
rect 240685 201456 240690 201512
rect 240746 201456 240874 201512
rect 240930 201456 240935 201512
rect 240685 201454 240935 201456
rect 240685 201451 240751 201454
rect 240869 201451 240935 201454
rect 264329 201514 264395 201517
rect 264513 201514 264579 201517
rect 264329 201512 264579 201514
rect 264329 201456 264334 201512
rect 264390 201456 264518 201512
rect 264574 201456 264579 201512
rect 264329 201454 264579 201456
rect 264329 201451 264395 201454
rect 264513 201451 264579 201454
rect 293125 201514 293191 201517
rect 293309 201514 293375 201517
rect 293125 201512 293375 201514
rect 293125 201456 293130 201512
rect 293186 201456 293314 201512
rect 293370 201456 293375 201512
rect 293125 201454 293375 201456
rect 293125 201451 293191 201454
rect 293309 201451 293375 201454
rect 294597 201514 294663 201517
rect 294781 201514 294847 201517
rect 294597 201512 294847 201514
rect 294597 201456 294602 201512
rect 294658 201456 294786 201512
rect 294842 201456 294847 201512
rect 294597 201454 294847 201456
rect 294597 201451 294663 201454
rect 294781 201451 294847 201454
rect 295885 201514 295951 201517
rect 296069 201514 296135 201517
rect 295885 201512 296135 201514
rect 295885 201456 295890 201512
rect 295946 201456 296074 201512
rect 296130 201456 296135 201512
rect 295885 201454 296135 201456
rect 320958 201514 321018 201590
rect 321093 201587 321159 201590
rect 321093 201514 321159 201517
rect 320958 201512 321159 201514
rect 320958 201456 321098 201512
rect 321154 201456 321159 201512
rect 320958 201454 321159 201456
rect 295885 201451 295951 201454
rect 296069 201451 296135 201454
rect 321093 201451 321159 201454
rect 322105 201514 322171 201517
rect 322289 201514 322355 201517
rect 322105 201512 322355 201514
rect 322105 201456 322110 201512
rect 322166 201456 322294 201512
rect 322350 201456 322355 201512
rect 322105 201454 322355 201456
rect 322105 201451 322171 201454
rect 322289 201451 322355 201454
rect 262857 200154 262923 200157
rect 263041 200154 263107 200157
rect 262857 200152 263107 200154
rect 262857 200096 262862 200152
rect 262918 200096 263046 200152
rect 263102 200096 263107 200152
rect 262857 200094 263107 200096
rect 262857 200091 262923 200094
rect 263041 200091 263107 200094
rect 301589 198794 301655 198797
rect 301773 198794 301839 198797
rect 301589 198792 301839 198794
rect 301589 198736 301594 198792
rect 301650 198736 301778 198792
rect 301834 198736 301839 198792
rect 301589 198734 301839 198736
rect 301589 198731 301655 198734
rect 301773 198731 301839 198734
rect -960 193898 480 193988
rect 2773 193898 2839 193901
rect -960 193896 2839 193898
rect -960 193840 2778 193896
rect 2834 193840 2839 193896
rect -960 193838 2839 193840
rect -960 193748 480 193838
rect 2773 193835 2839 193838
rect 583520 193476 584960 193716
rect 100661 193218 100727 193221
rect 100845 193218 100911 193221
rect 100661 193216 100911 193218
rect 100661 193160 100666 193216
rect 100722 193160 100850 193216
rect 100906 193160 100911 193216
rect 100661 193158 100911 193160
rect 100661 193155 100727 193158
rect 100845 193155 100911 193158
rect 244181 193218 244247 193221
rect 244457 193218 244523 193221
rect 244181 193216 244523 193218
rect 244181 193160 244186 193216
rect 244242 193160 244462 193216
rect 244518 193160 244523 193216
rect 244181 193158 244523 193160
rect 244181 193155 244247 193158
rect 244457 193155 244523 193158
rect 246389 193218 246455 193221
rect 246573 193218 246639 193221
rect 246389 193216 246639 193218
rect 246389 193160 246394 193216
rect 246450 193160 246578 193216
rect 246634 193160 246639 193216
rect 246389 193158 246639 193160
rect 246389 193155 246455 193158
rect 246573 193155 246639 193158
rect 294781 191994 294847 191997
rect 296069 191994 296135 191997
rect 294781 191992 294890 191994
rect 294781 191936 294786 191992
rect 294842 191936 294890 191992
rect 294781 191931 294890 191936
rect 296069 191992 296178 191994
rect 296069 191936 296074 191992
rect 296130 191936 296178 191992
rect 296069 191931 296178 191936
rect 294830 191861 294890 191931
rect 296118 191861 296178 191931
rect 107469 191858 107535 191861
rect 107653 191858 107719 191861
rect 107469 191856 107719 191858
rect 107469 191800 107474 191856
rect 107530 191800 107658 191856
rect 107714 191800 107719 191856
rect 107469 191798 107719 191800
rect 107469 191795 107535 191798
rect 107653 191795 107719 191798
rect 264329 191858 264395 191861
rect 264513 191858 264579 191861
rect 264329 191856 264579 191858
rect 264329 191800 264334 191856
rect 264390 191800 264518 191856
rect 264574 191800 264579 191856
rect 264329 191798 264579 191800
rect 264329 191795 264395 191798
rect 264513 191795 264579 191798
rect 293125 191858 293191 191861
rect 293309 191858 293375 191861
rect 293125 191856 293375 191858
rect 293125 191800 293130 191856
rect 293186 191800 293314 191856
rect 293370 191800 293375 191856
rect 293125 191798 293375 191800
rect 293125 191795 293191 191798
rect 293309 191795 293375 191798
rect 294781 191856 294890 191861
rect 294781 191800 294786 191856
rect 294842 191800 294890 191856
rect 294781 191798 294890 191800
rect 296069 191856 296178 191861
rect 296069 191800 296074 191856
rect 296130 191800 296178 191856
rect 296069 191798 296178 191800
rect 345381 191858 345447 191861
rect 345565 191858 345631 191861
rect 345381 191856 345631 191858
rect 345381 191800 345386 191856
rect 345442 191800 345570 191856
rect 345626 191800 345631 191856
rect 345381 191798 345631 191800
rect 294781 191795 294847 191798
rect 296069 191795 296135 191798
rect 345381 191795 345447 191798
rect 345565 191795 345631 191798
rect 335905 190498 335971 190501
rect 336089 190498 336155 190501
rect 335905 190496 336155 190498
rect 335905 190440 335910 190496
rect 335966 190440 336094 190496
rect 336150 190440 336155 190496
rect 335905 190438 336155 190440
rect 335905 190435 335971 190438
rect 336089 190435 336155 190438
rect 231209 183562 231275 183565
rect 231393 183562 231459 183565
rect 231209 183560 231459 183562
rect 231209 183504 231214 183560
rect 231270 183504 231398 183560
rect 231454 183504 231459 183560
rect 231209 183502 231459 183504
rect 231209 183499 231275 183502
rect 231393 183499 231459 183502
rect 245837 183562 245903 183565
rect 246021 183562 246087 183565
rect 245837 183560 246087 183562
rect 245837 183504 245842 183560
rect 245898 183504 246026 183560
rect 246082 183504 246087 183560
rect 245837 183502 246087 183504
rect 245837 183499 245903 183502
rect 246021 183499 246087 183502
rect 321093 182338 321159 182341
rect 320958 182336 321159 182338
rect 320958 182280 321098 182336
rect 321154 182280 321159 182336
rect 320958 182278 321159 182280
rect 232129 182202 232195 182205
rect 232313 182202 232379 182205
rect 232129 182200 232379 182202
rect 232129 182144 232134 182200
rect 232190 182144 232318 182200
rect 232374 182144 232379 182200
rect 232129 182142 232379 182144
rect 232129 182139 232195 182142
rect 232313 182139 232379 182142
rect 240685 182202 240751 182205
rect 240869 182202 240935 182205
rect 240685 182200 240935 182202
rect 240685 182144 240690 182200
rect 240746 182144 240874 182200
rect 240930 182144 240935 182200
rect 240685 182142 240935 182144
rect 240685 182139 240751 182142
rect 240869 182139 240935 182142
rect 264329 182202 264395 182205
rect 264513 182202 264579 182205
rect 264329 182200 264579 182202
rect 264329 182144 264334 182200
rect 264390 182144 264518 182200
rect 264574 182144 264579 182200
rect 264329 182142 264579 182144
rect 264329 182139 264395 182142
rect 264513 182139 264579 182142
rect 265617 182202 265683 182205
rect 265801 182202 265867 182205
rect 265617 182200 265867 182202
rect 265617 182144 265622 182200
rect 265678 182144 265806 182200
rect 265862 182144 265867 182200
rect 265617 182142 265867 182144
rect 265617 182139 265683 182142
rect 265801 182139 265867 182142
rect 293125 182202 293191 182205
rect 293309 182202 293375 182205
rect 293125 182200 293375 182202
rect 293125 182144 293130 182200
rect 293186 182144 293314 182200
rect 293370 182144 293375 182200
rect 293125 182142 293375 182144
rect 293125 182139 293191 182142
rect 293309 182139 293375 182142
rect 294597 182202 294663 182205
rect 294781 182202 294847 182205
rect 294597 182200 294847 182202
rect 294597 182144 294602 182200
rect 294658 182144 294786 182200
rect 294842 182144 294847 182200
rect 294597 182142 294847 182144
rect 294597 182139 294663 182142
rect 294781 182139 294847 182142
rect 295885 182202 295951 182205
rect 296069 182202 296135 182205
rect 295885 182200 296135 182202
rect 295885 182144 295890 182200
rect 295946 182144 296074 182200
rect 296130 182144 296135 182200
rect 295885 182142 296135 182144
rect 320958 182202 321018 182278
rect 321093 182275 321159 182278
rect 321093 182202 321159 182205
rect 320958 182200 321159 182202
rect 320958 182144 321098 182200
rect 321154 182144 321159 182200
rect 320958 182142 321159 182144
rect 295885 182139 295951 182142
rect 296069 182139 296135 182142
rect 321093 182139 321159 182142
rect 580625 181930 580691 181933
rect 583520 181930 584960 182020
rect 580625 181928 584960 181930
rect 580625 181872 580630 181928
rect 580686 181872 584960 181928
rect 580625 181870 584960 181872
rect 580625 181867 580691 181870
rect 583520 181780 584960 181870
rect -960 179482 480 179572
rect 2773 179482 2839 179485
rect -960 179480 2839 179482
rect -960 179424 2778 179480
rect 2834 179424 2839 179480
rect -960 179422 2839 179424
rect -960 179332 480 179422
rect 2773 179419 2839 179422
rect 100661 173906 100727 173909
rect 100845 173906 100911 173909
rect 100661 173904 100911 173906
rect 100661 173848 100666 173904
rect 100722 173848 100850 173904
rect 100906 173848 100911 173904
rect 100661 173846 100911 173848
rect 100661 173843 100727 173846
rect 100845 173843 100911 173846
rect 244181 173906 244247 173909
rect 244457 173906 244523 173909
rect 244181 173904 244523 173906
rect 244181 173848 244186 173904
rect 244242 173848 244462 173904
rect 244518 173848 244523 173904
rect 244181 173846 244523 173848
rect 244181 173843 244247 173846
rect 244457 173843 244523 173846
rect 107469 172546 107535 172549
rect 107653 172546 107719 172549
rect 107469 172544 107719 172546
rect 107469 172488 107474 172544
rect 107530 172488 107658 172544
rect 107714 172488 107719 172544
rect 107469 172486 107719 172488
rect 107469 172483 107535 172486
rect 107653 172483 107719 172486
rect 231945 172546 232011 172549
rect 232129 172546 232195 172549
rect 231945 172544 232195 172546
rect 231945 172488 231950 172544
rect 232006 172488 232134 172544
rect 232190 172488 232195 172544
rect 231945 172486 232195 172488
rect 231945 172483 232011 172486
rect 232129 172483 232195 172486
rect 371877 170234 371943 170237
rect 367142 170232 371943 170234
rect 367142 170176 371882 170232
rect 371938 170176 371943 170232
rect 367142 170174 371943 170176
rect 342662 169900 342668 169964
rect 342732 169962 342738 169964
rect 350441 169962 350507 169965
rect 342732 169960 350507 169962
rect 342732 169904 350446 169960
rect 350502 169904 350507 169960
rect 342732 169902 350507 169904
rect 342732 169900 342738 169902
rect 350441 169899 350507 169902
rect 367001 169962 367067 169965
rect 367142 169962 367202 170174
rect 371877 170171 371943 170174
rect 376702 170036 376708 170100
rect 376772 170098 376778 170100
rect 583520 170098 584960 170188
rect 376772 170038 393330 170098
rect 376772 170036 376778 170038
rect 367001 169960 367202 169962
rect 367001 169904 367006 169960
rect 367062 169904 367202 169960
rect 367001 169902 367202 169904
rect 393270 169962 393330 170038
rect 403022 170038 412650 170098
rect 393270 169902 402898 169962
rect 367001 169899 367067 169902
rect 350625 169826 350691 169829
rect 357382 169826 357388 169828
rect 350625 169824 357388 169826
rect 350625 169768 350630 169824
rect 350686 169768 357388 169824
rect 350625 169766 357388 169768
rect 350625 169763 350691 169766
rect 357382 169764 357388 169766
rect 357452 169764 357458 169828
rect 371877 169826 371943 169829
rect 376702 169826 376708 169828
rect 371877 169824 376708 169826
rect 371877 169768 371882 169824
rect 371938 169768 376708 169824
rect 371877 169766 376708 169768
rect 371877 169763 371943 169766
rect 376702 169764 376708 169766
rect 376772 169764 376778 169828
rect 402838 169826 402898 169902
rect 403022 169826 403082 170038
rect 412590 169962 412650 170038
rect 422342 170038 431970 170098
rect 412590 169902 422218 169962
rect 402838 169766 403082 169826
rect 422158 169826 422218 169902
rect 422342 169826 422402 170038
rect 431910 169962 431970 170038
rect 441662 170038 451290 170098
rect 431910 169902 441538 169962
rect 422158 169766 422402 169826
rect 441478 169826 441538 169902
rect 441662 169826 441722 170038
rect 451230 169962 451290 170038
rect 460982 170038 470610 170098
rect 451230 169902 460858 169962
rect 441478 169766 441722 169826
rect 460798 169826 460858 169902
rect 460982 169826 461042 170038
rect 470550 169962 470610 170038
rect 480302 170038 489930 170098
rect 470550 169902 480178 169962
rect 460798 169766 461042 169826
rect 480118 169826 480178 169902
rect 480302 169826 480362 170038
rect 489870 169962 489930 170038
rect 499622 170038 509250 170098
rect 489870 169902 499498 169962
rect 480118 169766 480362 169826
rect 499438 169826 499498 169902
rect 499622 169826 499682 170038
rect 509190 169962 509250 170038
rect 518942 170038 528570 170098
rect 509190 169902 518818 169962
rect 499438 169766 499682 169826
rect 518758 169826 518818 169902
rect 518942 169826 519002 170038
rect 528510 169962 528570 170038
rect 538262 170038 547890 170098
rect 528510 169902 538138 169962
rect 518758 169766 519002 169826
rect 538078 169826 538138 169902
rect 538262 169826 538322 170038
rect 547830 169962 547890 170038
rect 557582 170038 567210 170098
rect 547830 169902 557458 169962
rect 538078 169766 538322 169826
rect 557398 169826 557458 169902
rect 557582 169826 557642 170038
rect 567150 169962 567210 170038
rect 583342 170038 584960 170098
rect 583342 169962 583402 170038
rect 567150 169902 576778 169962
rect 557398 169766 557642 169826
rect 576718 169826 576778 169902
rect 576902 169902 583402 169962
rect 583520 169948 584960 170038
rect 576902 169826 576962 169902
rect 576718 169766 576962 169826
rect 357382 169492 357388 169556
rect 357452 169554 357458 169556
rect 367001 169554 367067 169557
rect 357452 169552 367067 169554
rect 357452 169496 367006 169552
rect 367062 169496 367067 169552
rect 357452 169494 367067 169496
rect 357452 169492 357458 169494
rect 367001 169491 367067 169494
rect -960 165066 480 165156
rect 3693 165066 3759 165069
rect -960 165064 3759 165066
rect -960 165008 3698 165064
rect 3754 165008 3759 165064
rect -960 165006 3759 165008
rect -960 164916 480 165006
rect 3693 165003 3759 165006
rect 244917 164386 244983 164389
rect 254761 164386 254827 164389
rect 258809 164386 258875 164389
rect 244917 164384 245026 164386
rect 244917 164328 244922 164384
rect 244978 164328 245026 164384
rect 244917 164323 245026 164328
rect 244966 164253 245026 164323
rect 254718 164384 254827 164386
rect 254718 164328 254766 164384
rect 254822 164328 254827 164384
rect 254718 164323 254827 164328
rect 258766 164384 258875 164386
rect 258766 164328 258814 164384
rect 258870 164328 258875 164384
rect 258766 164323 258875 164328
rect 254718 164253 254778 164323
rect 258766 164253 258826 164323
rect 100661 164250 100727 164253
rect 100845 164250 100911 164253
rect 100661 164248 100911 164250
rect 100661 164192 100666 164248
rect 100722 164192 100850 164248
rect 100906 164192 100911 164248
rect 100661 164190 100911 164192
rect 100661 164187 100727 164190
rect 100845 164187 100911 164190
rect 244181 164250 244247 164253
rect 244365 164250 244431 164253
rect 244181 164248 244431 164250
rect 244181 164192 244186 164248
rect 244242 164192 244370 164248
rect 244426 164192 244431 164248
rect 244181 164190 244431 164192
rect 244966 164248 245075 164253
rect 244966 164192 245014 164248
rect 245070 164192 245075 164248
rect 244966 164190 245075 164192
rect 254718 164248 254827 164253
rect 254718 164192 254766 164248
rect 254822 164192 254827 164248
rect 254718 164190 254827 164192
rect 258766 164248 258875 164253
rect 258766 164192 258814 164248
rect 258870 164192 258875 164248
rect 258766 164190 258875 164192
rect 244181 164187 244247 164190
rect 244365 164187 244431 164190
rect 245009 164187 245075 164190
rect 254761 164187 254827 164190
rect 258809 164187 258875 164190
rect 340137 164250 340203 164253
rect 340321 164250 340387 164253
rect 340137 164248 340387 164250
rect 340137 164192 340142 164248
rect 340198 164192 340326 164248
rect 340382 164192 340387 164248
rect 340137 164190 340387 164192
rect 340137 164187 340203 164190
rect 340321 164187 340387 164190
rect 240685 162890 240751 162893
rect 240869 162890 240935 162893
rect 240685 162888 240935 162890
rect 240685 162832 240690 162888
rect 240746 162832 240874 162888
rect 240930 162832 240935 162888
rect 240685 162830 240935 162832
rect 240685 162827 240751 162830
rect 240869 162827 240935 162830
rect 335905 161530 335971 161533
rect 336089 161530 336155 161533
rect 335905 161528 336155 161530
rect 335905 161472 335910 161528
rect 335966 161472 336094 161528
rect 336150 161472 336155 161528
rect 335905 161470 336155 161472
rect 335905 161467 335971 161470
rect 336089 161467 336155 161470
rect 322289 161394 322355 161397
rect 322289 161392 322490 161394
rect 322289 161336 322294 161392
rect 322350 161336 322490 161392
rect 322289 161334 322490 161336
rect 322289 161331 322355 161334
rect 322430 161261 322490 161334
rect 322381 161256 322490 161261
rect 322381 161200 322386 161256
rect 322442 161200 322490 161256
rect 322381 161198 322490 161200
rect 322381 161195 322447 161198
rect 580533 158402 580599 158405
rect 583520 158402 584960 158492
rect 580533 158400 584960 158402
rect 580533 158344 580538 158400
rect 580594 158344 584960 158400
rect 580533 158342 584960 158344
rect 580533 158339 580599 158342
rect 583520 158252 584960 158342
rect 246481 154730 246547 154733
rect 246438 154728 246547 154730
rect 246438 154672 246486 154728
rect 246542 154672 246547 154728
rect 246438 154667 246547 154672
rect 246438 154597 246498 154667
rect 244181 154594 244247 154597
rect 244457 154594 244523 154597
rect 244181 154592 244523 154594
rect 244181 154536 244186 154592
rect 244242 154536 244462 154592
rect 244518 154536 244523 154592
rect 244181 154534 244523 154536
rect 244181 154531 244247 154534
rect 244457 154531 244523 154534
rect 246389 154592 246498 154597
rect 246389 154536 246394 154592
rect 246450 154536 246498 154592
rect 246389 154534 246498 154536
rect 345381 154594 345447 154597
rect 345565 154594 345631 154597
rect 345381 154592 345631 154594
rect 345381 154536 345386 154592
rect 345442 154536 345570 154592
rect 345626 154536 345631 154592
rect 345381 154534 345631 154536
rect 246389 154531 246455 154534
rect 345381 154531 345447 154534
rect 345565 154531 345631 154534
rect -960 150786 480 150876
rect 2773 150786 2839 150789
rect -960 150784 2839 150786
rect -960 150728 2778 150784
rect 2834 150728 2839 150784
rect -960 150726 2839 150728
rect -960 150636 480 150726
rect 2773 150723 2839 150726
rect 583520 146556 584960 146796
rect 100661 144938 100727 144941
rect 100845 144938 100911 144941
rect 100661 144936 100911 144938
rect 100661 144880 100666 144936
rect 100722 144880 100850 144936
rect 100906 144880 100911 144936
rect 100661 144878 100911 144880
rect 100661 144875 100727 144878
rect 100845 144875 100911 144878
rect 231209 144938 231275 144941
rect 231393 144938 231459 144941
rect 231209 144936 231459 144938
rect 231209 144880 231214 144936
rect 231270 144880 231398 144936
rect 231454 144880 231459 144936
rect 231209 144878 231459 144880
rect 231209 144875 231275 144878
rect 231393 144875 231459 144878
rect 340137 144938 340203 144941
rect 340413 144938 340479 144941
rect 340137 144936 340479 144938
rect 340137 144880 340142 144936
rect 340198 144880 340418 144936
rect 340474 144880 340479 144936
rect 340137 144878 340479 144880
rect 340137 144875 340203 144878
rect 340413 144875 340479 144878
rect 319621 143714 319687 143717
rect 319621 143712 319730 143714
rect 319621 143656 319626 143712
rect 319682 143656 319730 143712
rect 319621 143651 319730 143656
rect 319670 143581 319730 143651
rect 240685 143578 240751 143581
rect 240869 143578 240935 143581
rect 240685 143576 240935 143578
rect 240685 143520 240690 143576
rect 240746 143520 240874 143576
rect 240930 143520 240935 143576
rect 240685 143518 240935 143520
rect 240685 143515 240751 143518
rect 240869 143515 240935 143518
rect 319621 143576 319730 143581
rect 319621 143520 319626 143576
rect 319682 143520 319730 143576
rect 319621 143518 319730 143520
rect 319621 143515 319687 143518
rect 320909 142218 320975 142221
rect 320909 142216 321018 142218
rect 320909 142160 320914 142216
rect 320970 142160 321018 142216
rect 320909 142155 321018 142160
rect 320958 141949 321018 142155
rect 320958 141944 321067 141949
rect 320958 141888 321006 141944
rect 321062 141888 321067 141944
rect 320958 141886 321067 141888
rect 321001 141883 321067 141886
rect 301957 141266 302023 141269
rect 301822 141264 302023 141266
rect 301822 141208 301962 141264
rect 302018 141208 302023 141264
rect 301822 141206 302023 141208
rect 301822 140858 301882 141206
rect 301957 141203 302023 141206
rect 301957 140858 302023 140861
rect 301822 140856 302023 140858
rect 301822 140800 301962 140856
rect 302018 140800 302023 140856
rect 301822 140798 302023 140800
rect 301957 140795 302023 140798
rect 232497 139634 232563 139637
rect 232454 139632 232563 139634
rect 232454 139576 232502 139632
rect 232558 139576 232563 139632
rect 232454 139571 232563 139576
rect 232454 139501 232514 139571
rect 232454 139496 232563 139501
rect 232454 139440 232502 139496
rect 232558 139440 232563 139496
rect 232454 139438 232563 139440
rect 232497 139435 232563 139438
rect 244457 138684 244523 138685
rect 244406 138620 244412 138684
rect 244476 138682 244523 138684
rect 244476 138680 244568 138682
rect 244518 138624 244568 138680
rect 244476 138622 244568 138624
rect 244476 138620 244523 138622
rect 244457 138619 244523 138620
rect 232589 136642 232655 136645
rect 232865 136642 232931 136645
rect 232589 136640 232931 136642
rect 232589 136584 232594 136640
rect 232650 136584 232870 136640
rect 232926 136584 232931 136640
rect 232589 136582 232931 136584
rect 232589 136579 232655 136582
rect 232865 136579 232931 136582
rect -960 136370 480 136460
rect 2773 136370 2839 136373
rect -960 136368 2839 136370
rect -960 136312 2778 136368
rect 2834 136312 2839 136368
rect -960 136310 2839 136312
rect -960 136220 480 136310
rect 2773 136307 2839 136310
rect 580441 134874 580507 134877
rect 583520 134874 584960 134964
rect 580441 134872 584960 134874
rect 580441 134816 580446 134872
rect 580502 134816 584960 134872
rect 580441 134814 584960 134816
rect 580441 134811 580507 134814
rect 583520 134724 584960 134814
rect 100661 125626 100727 125629
rect 100845 125626 100911 125629
rect 100661 125624 100911 125626
rect 100661 125568 100666 125624
rect 100722 125568 100850 125624
rect 100906 125568 100911 125624
rect 100661 125566 100911 125568
rect 100661 125563 100727 125566
rect 100845 125563 100911 125566
rect 231209 125626 231275 125629
rect 231393 125626 231459 125629
rect 244365 125628 244431 125629
rect 244365 125626 244412 125628
rect 231209 125624 231459 125626
rect 231209 125568 231214 125624
rect 231270 125568 231398 125624
rect 231454 125568 231459 125624
rect 231209 125566 231459 125568
rect 244320 125624 244412 125626
rect 244320 125568 244370 125624
rect 244320 125566 244412 125568
rect 231209 125563 231275 125566
rect 231393 125563 231459 125566
rect 244365 125564 244412 125566
rect 244476 125564 244482 125628
rect 244365 125563 244431 125564
rect 245837 124266 245903 124269
rect 246021 124266 246087 124269
rect 245837 124264 246087 124266
rect 245837 124208 245842 124264
rect 245898 124208 246026 124264
rect 246082 124208 246087 124264
rect 245837 124206 246087 124208
rect 245837 124203 245903 124206
rect 246021 124203 246087 124206
rect 256969 124266 257035 124269
rect 257153 124266 257219 124269
rect 256969 124264 257219 124266
rect 256969 124208 256974 124264
rect 257030 124208 257158 124264
rect 257214 124208 257219 124264
rect 256969 124206 257219 124208
rect 256969 124203 257035 124206
rect 257153 124203 257219 124206
rect 345289 124266 345355 124269
rect 345565 124266 345631 124269
rect 345289 124264 345631 124266
rect 345289 124208 345294 124264
rect 345350 124208 345570 124264
rect 345626 124208 345631 124264
rect 345289 124206 345631 124208
rect 345289 124203 345355 124206
rect 345565 124203 345631 124206
rect 579613 123178 579679 123181
rect 583520 123178 584960 123268
rect 579613 123176 584960 123178
rect 579613 123120 579618 123176
rect 579674 123120 584960 123176
rect 579613 123118 584960 123120
rect 579613 123115 579679 123118
rect 583520 123028 584960 123118
rect -960 122090 480 122180
rect 3601 122090 3667 122093
rect -960 122088 3667 122090
rect -960 122032 3606 122088
rect 3662 122032 3667 122088
rect -960 122030 3667 122032
rect -960 121940 480 122030
rect 3601 122027 3667 122030
rect 320909 113250 320975 113253
rect 321093 113250 321159 113253
rect 320909 113248 321159 113250
rect 320909 113192 320914 113248
rect 320970 113192 321098 113248
rect 321154 113192 321159 113248
rect 320909 113190 321159 113192
rect 320909 113187 320975 113190
rect 321093 113187 321159 113190
rect 580349 111482 580415 111485
rect 583520 111482 584960 111572
rect 580349 111480 584960 111482
rect 580349 111424 580354 111480
rect 580410 111424 584960 111480
rect 580349 111422 584960 111424
rect 580349 111419 580415 111422
rect 583520 111332 584960 111422
rect -960 107674 480 107764
rect 3325 107674 3391 107677
rect -960 107672 3391 107674
rect -960 107616 3330 107672
rect 3386 107616 3391 107672
rect -960 107614 3391 107616
rect -960 107524 480 107614
rect 3325 107611 3391 107614
rect 232681 107674 232747 107677
rect 232865 107674 232931 107677
rect 232681 107672 232931 107674
rect 232681 107616 232686 107672
rect 232742 107616 232870 107672
rect 232926 107616 232931 107672
rect 232681 107614 232931 107616
rect 232681 107611 232747 107614
rect 232865 107611 232931 107614
rect 583520 99636 584960 99876
rect 258717 93802 258783 93805
rect 258901 93802 258967 93805
rect 258717 93800 258967 93802
rect 258717 93744 258722 93800
rect 258778 93744 258906 93800
rect 258962 93744 258967 93800
rect 258717 93742 258967 93744
rect 258717 93739 258783 93742
rect 258901 93739 258967 93742
rect -960 93258 480 93348
rect 3509 93258 3575 93261
rect -960 93256 3575 93258
rect -960 93200 3514 93256
rect 3570 93200 3575 93256
rect -960 93198 3575 93200
rect -960 93108 480 93198
rect 3509 93195 3575 93198
rect 233734 90476 233740 90540
rect 233804 90538 233810 90540
rect 238661 90538 238727 90541
rect 233804 90536 238727 90538
rect 233804 90480 238666 90536
rect 238722 90480 238727 90536
rect 233804 90478 238727 90480
rect 233804 90476 233810 90478
rect 238661 90475 238727 90478
rect 583520 87954 584960 88044
rect 583342 87894 584960 87954
rect 365662 87348 365668 87412
rect 365732 87410 365738 87412
rect 375281 87410 375347 87413
rect 365732 87408 375347 87410
rect 365732 87352 375286 87408
rect 375342 87352 375347 87408
rect 365732 87350 375347 87352
rect 365732 87348 365738 87350
rect 375281 87347 375347 87350
rect 386321 87274 386387 87277
rect 386321 87272 393330 87274
rect 386321 87216 386326 87272
rect 386382 87216 393330 87272
rect 386321 87214 393330 87216
rect 386321 87211 386387 87214
rect 238661 87138 238727 87141
rect 350441 87138 350507 87141
rect 238661 87136 244842 87138
rect 238661 87080 238666 87136
rect 238722 87080 244842 87136
rect 238661 87078 244842 87080
rect 238661 87075 238727 87078
rect 244782 87002 244842 87078
rect 330526 87136 350507 87138
rect 330526 87080 350446 87136
rect 350502 87080 350507 87136
rect 330526 87078 350507 87080
rect 249701 87002 249767 87005
rect 244782 87000 249767 87002
rect 244782 86944 249706 87000
rect 249762 86944 249767 87000
rect 244782 86942 249767 86944
rect 249701 86939 249767 86942
rect 259453 87002 259519 87005
rect 330526 87002 330586 87078
rect 350441 87075 350507 87078
rect 360285 87138 360351 87141
rect 365662 87138 365668 87140
rect 360285 87136 365668 87138
rect 360285 87080 360290 87136
rect 360346 87080 365668 87136
rect 360285 87078 365668 87080
rect 360285 87075 360351 87078
rect 365662 87076 365668 87078
rect 365732 87076 365738 87140
rect 379421 87138 379487 87141
rect 376710 87136 379487 87138
rect 376710 87080 379426 87136
rect 379482 87080 379487 87136
rect 376710 87078 379487 87080
rect 393270 87138 393330 87214
rect 403022 87214 412650 87274
rect 393270 87078 402898 87138
rect 259453 87000 330586 87002
rect 259453 86944 259458 87000
rect 259514 86944 330586 87000
rect 259453 86942 330586 86944
rect 350625 87002 350691 87005
rect 360101 87002 360167 87005
rect 350625 87000 360167 87002
rect 350625 86944 350630 87000
rect 350686 86944 360106 87000
rect 360162 86944 360167 87000
rect 350625 86942 360167 86944
rect 259453 86939 259519 86942
rect 350625 86939 350691 86942
rect 360101 86939 360167 86942
rect 375281 87002 375347 87005
rect 376710 87002 376770 87078
rect 379421 87075 379487 87078
rect 375281 87000 376770 87002
rect 375281 86944 375286 87000
rect 375342 86944 376770 87000
rect 375281 86942 376770 86944
rect 402838 87002 402898 87078
rect 403022 87002 403082 87214
rect 412590 87138 412650 87214
rect 422342 87214 431970 87274
rect 412590 87078 422218 87138
rect 402838 86942 403082 87002
rect 422158 87002 422218 87078
rect 422342 87002 422402 87214
rect 431910 87138 431970 87214
rect 441662 87214 451290 87274
rect 431910 87078 441538 87138
rect 422158 86942 422402 87002
rect 441478 87002 441538 87078
rect 441662 87002 441722 87214
rect 451230 87138 451290 87214
rect 460982 87214 470610 87274
rect 451230 87078 460858 87138
rect 441478 86942 441722 87002
rect 460798 87002 460858 87078
rect 460982 87002 461042 87214
rect 470550 87138 470610 87214
rect 480302 87214 489930 87274
rect 470550 87078 480178 87138
rect 460798 86942 461042 87002
rect 480118 87002 480178 87078
rect 480302 87002 480362 87214
rect 489870 87138 489930 87214
rect 499622 87214 509250 87274
rect 489870 87078 499498 87138
rect 480118 86942 480362 87002
rect 499438 87002 499498 87078
rect 499622 87002 499682 87214
rect 509190 87138 509250 87214
rect 518942 87214 528570 87274
rect 509190 87078 518818 87138
rect 499438 86942 499682 87002
rect 518758 87002 518818 87078
rect 518942 87002 519002 87214
rect 528510 87138 528570 87214
rect 538262 87214 547890 87274
rect 528510 87078 538138 87138
rect 518758 86942 519002 87002
rect 538078 87002 538138 87078
rect 538262 87002 538322 87214
rect 547830 87138 547890 87214
rect 557582 87214 567210 87274
rect 547830 87078 557458 87138
rect 538078 86942 538322 87002
rect 557398 87002 557458 87078
rect 557582 87002 557642 87214
rect 567150 87138 567210 87214
rect 583342 87138 583402 87894
rect 583520 87804 584960 87894
rect 567150 87078 576778 87138
rect 557398 86942 557642 87002
rect 576718 87002 576778 87078
rect 576902 87078 583402 87138
rect 576902 87002 576962 87078
rect 576718 86942 576962 87002
rect 375281 86939 375347 86942
rect 252093 86866 252159 86869
rect 259453 86866 259519 86869
rect 252093 86864 259519 86866
rect 252093 86808 252098 86864
rect 252154 86808 259458 86864
rect 259514 86808 259519 86864
rect 252093 86806 259519 86808
rect 252093 86803 252159 86806
rect 259453 86803 259519 86806
rect 3509 80066 3575 80069
rect 343582 80066 343588 80068
rect 3509 80064 343588 80066
rect 3509 80008 3514 80064
rect 3570 80008 343588 80064
rect 3509 80006 343588 80008
rect 3509 80003 3575 80006
rect 343582 80004 343588 80006
rect 343652 80004 343658 80068
rect -960 78978 480 79068
rect 3509 78978 3575 78981
rect -960 78976 3575 78978
rect -960 78920 3514 78976
rect 3570 78920 3575 78976
rect -960 78918 3575 78920
rect -960 78828 480 78918
rect 3509 78915 3575 78918
rect 246389 77618 246455 77621
rect 246389 77616 246498 77618
rect 246389 77560 246394 77616
rect 246450 77560 246498 77616
rect 246389 77555 246498 77560
rect 246438 77349 246498 77555
rect 246389 77344 246498 77349
rect 246389 77288 246394 77344
rect 246450 77288 246498 77344
rect 246389 77286 246498 77288
rect 246389 77283 246455 77286
rect 580257 76258 580323 76261
rect 583520 76258 584960 76348
rect 580257 76256 584960 76258
rect 580257 76200 580262 76256
rect 580318 76200 584960 76256
rect 580257 76198 584960 76200
rect 580257 76195 580323 76198
rect 583520 76108 584960 76198
rect 265801 74626 265867 74629
rect 266353 74626 266419 74629
rect 265801 74624 266419 74626
rect 265801 74568 265806 74624
rect 265862 74568 266358 74624
rect 266414 74568 266419 74624
rect 265801 74566 266419 74568
rect 265801 74563 265867 74566
rect 266353 74563 266419 74566
rect 265617 64970 265683 64973
rect 265801 64970 265867 64973
rect 265617 64968 265867 64970
rect 265617 64912 265622 64968
rect 265678 64912 265806 64968
rect 265862 64912 265867 64968
rect 265617 64910 265867 64912
rect 265617 64907 265683 64910
rect 265801 64907 265867 64910
rect 345238 64834 345244 64836
rect 614 64774 345244 64834
rect -960 64562 480 64652
rect 614 64562 674 64774
rect 345238 64772 345244 64774
rect 345308 64772 345314 64836
rect 583520 64562 584960 64652
rect -960 64502 674 64562
rect 583342 64502 584960 64562
rect -960 64412 480 64502
rect 324262 63956 324268 64020
rect 324332 64018 324338 64020
rect 333881 64018 333947 64021
rect 324332 64016 333947 64018
rect 324332 63960 333886 64016
rect 333942 63960 333947 64016
rect 324332 63958 333947 63960
rect 324332 63956 324338 63958
rect 333881 63955 333947 63958
rect 343582 63956 343588 64020
rect 343652 64018 343658 64020
rect 353201 64018 353267 64021
rect 371877 64018 371943 64021
rect 343652 64016 353267 64018
rect 343652 63960 353206 64016
rect 353262 63960 353267 64016
rect 343652 63958 353267 63960
rect 343652 63956 343658 63958
rect 353201 63955 353267 63958
rect 367142 64016 371943 64018
rect 367142 63960 371882 64016
rect 371938 63960 371943 64016
rect 367142 63958 371943 63960
rect 233918 63684 233924 63748
rect 233988 63746 233994 63748
rect 258022 63746 258028 63748
rect 233988 63686 258028 63746
rect 233988 63684 233994 63686
rect 258022 63684 258028 63686
rect 258092 63684 258098 63748
rect 278865 63746 278931 63749
rect 278822 63744 278931 63746
rect 278822 63688 278870 63744
rect 278926 63688 278931 63744
rect 278822 63683 278931 63688
rect 315982 63684 315988 63748
rect 316052 63746 316058 63748
rect 324262 63746 324268 63748
rect 316052 63686 324268 63746
rect 316052 63684 316058 63686
rect 324262 63684 324268 63686
rect 324332 63684 324338 63748
rect 333881 63746 333947 63749
rect 343582 63746 343588 63748
rect 333881 63744 343588 63746
rect 333881 63688 333886 63744
rect 333942 63688 343588 63744
rect 333881 63686 343588 63688
rect 333881 63683 333947 63686
rect 343582 63684 343588 63686
rect 343652 63684 343658 63748
rect 353201 63746 353267 63749
rect 354581 63746 354647 63749
rect 353201 63744 354647 63746
rect 353201 63688 353206 63744
rect 353262 63688 354586 63744
rect 354642 63688 354647 63744
rect 353201 63686 354647 63688
rect 353201 63683 353267 63686
rect 354581 63683 354647 63686
rect 367001 63746 367067 63749
rect 367142 63746 367202 63958
rect 371877 63955 371943 63958
rect 376702 63820 376708 63884
rect 376772 63882 376778 63884
rect 376772 63822 393330 63882
rect 376772 63820 376778 63822
rect 367001 63744 367202 63746
rect 367001 63688 367006 63744
rect 367062 63688 367202 63744
rect 367001 63686 367202 63688
rect 393270 63746 393330 63822
rect 403022 63822 412650 63882
rect 393270 63686 402898 63746
rect 367001 63683 367067 63686
rect 267733 63610 267799 63613
rect 267598 63608 267799 63610
rect 267598 63552 267738 63608
rect 267794 63552 267799 63608
rect 267598 63550 267799 63552
rect 258022 63412 258028 63476
rect 258092 63474 258098 63476
rect 267598 63474 267658 63550
rect 267733 63547 267799 63550
rect 277158 63548 277164 63612
rect 277228 63610 277234 63612
rect 278822 63610 278882 63683
rect 277228 63550 278882 63610
rect 278957 63610 279023 63613
rect 354581 63610 354647 63613
rect 371877 63610 371943 63613
rect 376702 63610 376708 63612
rect 278957 63608 307770 63610
rect 278957 63552 278962 63608
rect 279018 63552 307770 63608
rect 278957 63550 307770 63552
rect 277228 63548 277234 63550
rect 278957 63547 279023 63550
rect 258092 63414 267658 63474
rect 258092 63412 258098 63414
rect 307710 63338 307770 63550
rect 354581 63608 354690 63610
rect 354581 63552 354586 63608
rect 354642 63552 354690 63608
rect 354581 63547 354690 63552
rect 371877 63608 376708 63610
rect 371877 63552 371882 63608
rect 371938 63552 376708 63608
rect 371877 63550 376708 63552
rect 371877 63547 371943 63550
rect 376702 63548 376708 63550
rect 376772 63548 376778 63612
rect 402838 63610 402898 63686
rect 403022 63610 403082 63822
rect 412590 63746 412650 63822
rect 422342 63822 431970 63882
rect 412590 63686 422218 63746
rect 402838 63550 403082 63610
rect 422158 63610 422218 63686
rect 422342 63610 422402 63822
rect 431910 63746 431970 63822
rect 441662 63822 451290 63882
rect 431910 63686 441538 63746
rect 422158 63550 422402 63610
rect 441478 63610 441538 63686
rect 441662 63610 441722 63822
rect 451230 63746 451290 63822
rect 460982 63822 470610 63882
rect 451230 63686 460858 63746
rect 441478 63550 441722 63610
rect 460798 63610 460858 63686
rect 460982 63610 461042 63822
rect 470550 63746 470610 63822
rect 480302 63822 489930 63882
rect 470550 63686 480178 63746
rect 460798 63550 461042 63610
rect 480118 63610 480178 63686
rect 480302 63610 480362 63822
rect 489870 63746 489930 63822
rect 499622 63822 509250 63882
rect 489870 63686 499498 63746
rect 480118 63550 480362 63610
rect 499438 63610 499498 63686
rect 499622 63610 499682 63822
rect 509190 63746 509250 63822
rect 518942 63822 528570 63882
rect 509190 63686 518818 63746
rect 499438 63550 499682 63610
rect 518758 63610 518818 63686
rect 518942 63610 519002 63822
rect 528510 63746 528570 63822
rect 538262 63822 547890 63882
rect 528510 63686 538138 63746
rect 518758 63550 519002 63610
rect 538078 63610 538138 63686
rect 538262 63610 538322 63822
rect 547830 63746 547890 63822
rect 557582 63822 567210 63882
rect 547830 63686 557458 63746
rect 538078 63550 538322 63610
rect 557398 63610 557458 63686
rect 557582 63610 557642 63822
rect 567150 63746 567210 63822
rect 583342 63746 583402 64502
rect 583520 64412 584960 64502
rect 567150 63686 576778 63746
rect 557398 63550 557642 63610
rect 576718 63610 576778 63686
rect 576902 63686 583402 63746
rect 576902 63610 576962 63686
rect 576718 63550 576962 63610
rect 354630 63474 354690 63547
rect 364241 63474 364307 63477
rect 354630 63472 364307 63474
rect 354630 63416 364246 63472
rect 364302 63416 364307 63472
rect 354630 63414 364307 63416
rect 364241 63411 364307 63414
rect 315982 63338 315988 63340
rect 307710 63278 315988 63338
rect 315982 63276 315988 63278
rect 316052 63276 316058 63340
rect 364241 63338 364307 63341
rect 367001 63338 367067 63341
rect 364241 63336 367067 63338
rect 364241 63280 364246 63336
rect 364302 63280 367006 63336
rect 367062 63280 367067 63336
rect 364241 63278 367067 63280
rect 364241 63275 364307 63278
rect 367001 63275 367067 63278
rect 267733 63202 267799 63205
rect 277158 63202 277164 63204
rect 267733 63200 277164 63202
rect 267733 63144 267738 63200
rect 267794 63144 277164 63200
rect 267733 63142 277164 63144
rect 267733 63139 267799 63142
rect 277158 63140 277164 63142
rect 277228 63140 277234 63204
rect 329005 62114 329071 62117
rect 329189 62114 329255 62117
rect 329005 62112 329255 62114
rect 329005 62056 329010 62112
rect 329066 62056 329194 62112
rect 329250 62056 329255 62112
rect 329005 62054 329255 62056
rect 329005 62051 329071 62054
rect 329189 62051 329255 62054
rect 583520 52716 584960 52956
rect 3325 50962 3391 50965
rect 345422 50962 345428 50964
rect 3325 50960 345428 50962
rect 3325 50904 3330 50960
rect 3386 50904 345428 50960
rect 3325 50902 345428 50904
rect 3325 50899 3391 50902
rect 345422 50900 345428 50902
rect 345492 50900 345498 50964
rect -960 50146 480 50236
rect 3325 50146 3391 50149
rect -960 50144 3391 50146
rect -960 50088 3330 50144
rect 3386 50088 3391 50144
rect -960 50086 3391 50088
rect -960 49996 480 50086
rect 3325 50083 3391 50086
rect 583520 41034 584960 41124
rect 583342 40974 584960 41034
rect 256601 40626 256667 40629
rect 355961 40626 356027 40629
rect 246990 40624 256667 40626
rect 246990 40568 256606 40624
rect 256662 40568 256667 40624
rect 246990 40566 256667 40568
rect 246990 40493 247050 40566
rect 256601 40563 256667 40566
rect 346350 40624 356027 40626
rect 346350 40568 355966 40624
rect 356022 40568 356027 40624
rect 346350 40566 356027 40568
rect 237414 40428 237420 40492
rect 237484 40490 237490 40492
rect 246941 40490 247050 40493
rect 237484 40488 247050 40490
rect 237484 40432 246946 40488
rect 247002 40432 247050 40488
rect 237484 40430 247050 40432
rect 237484 40428 237490 40430
rect 246941 40427 247050 40430
rect 267733 40490 267799 40493
rect 277158 40490 277164 40492
rect 267733 40488 277164 40490
rect 267733 40432 267738 40488
rect 267794 40432 277164 40488
rect 267733 40430 277164 40432
rect 267733 40427 267799 40430
rect 277158 40428 277164 40430
rect 277228 40428 277234 40492
rect 246990 40357 247050 40427
rect 246941 40354 247050 40357
rect 333881 40354 333947 40357
rect 246860 40352 247050 40354
rect 246860 40296 246946 40352
rect 247002 40296 247050 40352
rect 246860 40294 247050 40296
rect 307710 40352 333947 40354
rect 307710 40296 333886 40352
rect 333942 40296 333947 40352
rect 307710 40294 333947 40296
rect 246941 40291 247007 40294
rect 256601 40218 256667 40221
rect 259453 40218 259519 40221
rect 256601 40216 259519 40218
rect 256601 40160 256606 40216
rect 256662 40160 259458 40216
rect 259514 40160 259519 40216
rect 256601 40158 259519 40160
rect 256601 40155 256667 40158
rect 259453 40155 259519 40158
rect 283557 40218 283623 40221
rect 287053 40218 287119 40221
rect 283557 40216 287119 40218
rect 283557 40160 283562 40216
rect 283618 40160 287058 40216
rect 287114 40160 287119 40216
rect 283557 40158 287119 40160
rect 283557 40155 283623 40158
rect 287053 40155 287119 40158
rect 259453 40082 259519 40085
rect 267733 40082 267799 40085
rect 259453 40080 267799 40082
rect 259453 40024 259458 40080
rect 259514 40024 267738 40080
rect 267794 40024 267799 40080
rect 259453 40022 267799 40024
rect 259453 40019 259519 40022
rect 267733 40019 267799 40022
rect 277158 40020 277164 40084
rect 277228 40082 277234 40084
rect 307710 40082 307770 40294
rect 333881 40291 333947 40294
rect 344921 40354 344987 40357
rect 346350 40354 346410 40566
rect 355961 40563 356027 40566
rect 371877 40490 371943 40493
rect 344921 40352 346410 40354
rect 344921 40296 344926 40352
rect 344982 40296 346410 40352
rect 344921 40294 346410 40296
rect 367142 40488 371943 40490
rect 367142 40432 371882 40488
rect 371938 40432 371943 40488
rect 367142 40430 371943 40432
rect 344921 40291 344987 40294
rect 333881 40218 333947 40221
rect 335445 40218 335511 40221
rect 333881 40216 335511 40218
rect 333881 40160 333886 40216
rect 333942 40160 335450 40216
rect 335506 40160 335511 40216
rect 333881 40158 335511 40160
rect 333881 40155 333947 40158
rect 335445 40155 335511 40158
rect 367001 40218 367067 40221
rect 367142 40218 367202 40430
rect 371877 40427 371943 40430
rect 376702 40292 376708 40356
rect 376772 40354 376778 40356
rect 376772 40294 393330 40354
rect 376772 40292 376778 40294
rect 367001 40216 367202 40218
rect 367001 40160 367006 40216
rect 367062 40160 367202 40216
rect 367001 40158 367202 40160
rect 393270 40218 393330 40294
rect 403022 40294 412650 40354
rect 393270 40158 402898 40218
rect 367001 40155 367067 40158
rect 277228 40022 278882 40082
rect 277228 40020 277234 40022
rect 231710 39884 231716 39948
rect 231780 39946 231786 39948
rect 237414 39946 237420 39948
rect 231780 39886 237420 39946
rect 231780 39884 231786 39886
rect 237414 39884 237420 39886
rect 237484 39884 237490 39948
rect 278822 39810 278882 40022
rect 296486 40022 307770 40082
rect 355961 40082 356027 40085
rect 357382 40082 357388 40084
rect 355961 40080 357388 40082
rect 355961 40024 355966 40080
rect 356022 40024 357388 40080
rect 355961 40022 357388 40024
rect 283557 39810 283623 39813
rect 278822 39808 283623 39810
rect 278822 39752 283562 39808
rect 283618 39752 283623 39808
rect 278822 39750 283623 39752
rect 283557 39747 283623 39750
rect 287053 39674 287119 39677
rect 296486 39674 296546 40022
rect 355961 40019 356027 40022
rect 357382 40020 357388 40022
rect 357452 40020 357458 40084
rect 371877 40082 371943 40085
rect 376702 40082 376708 40084
rect 371877 40080 376708 40082
rect 371877 40024 371882 40080
rect 371938 40024 376708 40080
rect 371877 40022 376708 40024
rect 371877 40019 371943 40022
rect 376702 40020 376708 40022
rect 376772 40020 376778 40084
rect 402838 40082 402898 40158
rect 403022 40082 403082 40294
rect 412590 40218 412650 40294
rect 422342 40294 431970 40354
rect 412590 40158 422218 40218
rect 402838 40022 403082 40082
rect 422158 40082 422218 40158
rect 422342 40082 422402 40294
rect 431910 40218 431970 40294
rect 441662 40294 451290 40354
rect 431910 40158 441538 40218
rect 422158 40022 422402 40082
rect 441478 40082 441538 40158
rect 441662 40082 441722 40294
rect 451230 40218 451290 40294
rect 460982 40294 470610 40354
rect 451230 40158 460858 40218
rect 441478 40022 441722 40082
rect 460798 40082 460858 40158
rect 460982 40082 461042 40294
rect 470550 40218 470610 40294
rect 480302 40294 489930 40354
rect 470550 40158 480178 40218
rect 460798 40022 461042 40082
rect 480118 40082 480178 40158
rect 480302 40082 480362 40294
rect 489870 40218 489930 40294
rect 499622 40294 509250 40354
rect 489870 40158 499498 40218
rect 480118 40022 480362 40082
rect 499438 40082 499498 40158
rect 499622 40082 499682 40294
rect 509190 40218 509250 40294
rect 518942 40294 528570 40354
rect 509190 40158 518818 40218
rect 499438 40022 499682 40082
rect 518758 40082 518818 40158
rect 518942 40082 519002 40294
rect 528510 40218 528570 40294
rect 538262 40294 547890 40354
rect 528510 40158 538138 40218
rect 518758 40022 519002 40082
rect 538078 40082 538138 40158
rect 538262 40082 538322 40294
rect 547830 40218 547890 40294
rect 557582 40294 567210 40354
rect 547830 40158 557458 40218
rect 538078 40022 538322 40082
rect 557398 40082 557458 40158
rect 557582 40082 557642 40294
rect 567150 40218 567210 40294
rect 583342 40218 583402 40974
rect 583520 40884 584960 40974
rect 567150 40158 576778 40218
rect 557398 40022 557642 40082
rect 576718 40082 576778 40158
rect 576902 40158 583402 40218
rect 576902 40082 576962 40158
rect 576718 40022 576962 40082
rect 357382 39748 357388 39812
rect 357452 39810 357458 39812
rect 367001 39810 367067 39813
rect 357452 39808 367067 39810
rect 357452 39752 367006 39808
rect 367062 39752 367067 39808
rect 357452 39750 367067 39752
rect 357452 39748 357458 39750
rect 367001 39747 367067 39750
rect 287053 39672 296546 39674
rect 287053 39616 287058 39672
rect 287114 39616 296546 39672
rect 287053 39614 296546 39616
rect 287053 39611 287119 39614
rect -960 35866 480 35956
rect 347078 35866 347084 35868
rect -960 35806 347084 35866
rect -960 35716 480 35806
rect 347078 35804 347084 35806
rect 347148 35804 347154 35868
rect 329189 34506 329255 34509
rect 329373 34506 329439 34509
rect 329189 34504 329439 34506
rect 329189 34448 329194 34504
rect 329250 34448 329378 34504
rect 329434 34448 329439 34504
rect 329189 34446 329439 34448
rect 329189 34443 329255 34446
rect 329373 34443 329439 34446
rect 241462 29412 241468 29476
rect 241532 29474 241538 29476
rect 254485 29474 254551 29477
rect 355961 29474 356027 29477
rect 241532 29472 254551 29474
rect 241532 29416 254490 29472
rect 254546 29416 254551 29472
rect 241532 29414 254551 29416
rect 241532 29412 241538 29414
rect 254485 29411 254551 29414
rect 322062 29414 330586 29474
rect 232998 29140 233004 29204
rect 233068 29202 233074 29204
rect 241462 29202 241468 29204
rect 233068 29142 241468 29202
rect 233068 29140 233074 29142
rect 241462 29140 241468 29142
rect 241532 29140 241538 29204
rect 254485 29066 254551 29069
rect 322062 29066 322122 29414
rect 330526 29338 330586 29414
rect 346350 29472 356027 29474
rect 346350 29416 355966 29472
rect 356022 29416 356027 29472
rect 346350 29414 356027 29416
rect 337929 29338 337995 29341
rect 330526 29336 337995 29338
rect 330526 29280 337934 29336
rect 337990 29280 337995 29336
rect 330526 29278 337995 29280
rect 337929 29275 337995 29278
rect 338113 29338 338179 29341
rect 338113 29336 341626 29338
rect 338113 29280 338118 29336
rect 338174 29280 341626 29336
rect 338113 29278 341626 29280
rect 338113 29275 338179 29278
rect 341566 29202 341626 29278
rect 346350 29202 346410 29414
rect 355961 29411 356027 29414
rect 365662 29412 365668 29476
rect 365732 29474 365738 29476
rect 375281 29474 375347 29477
rect 365732 29472 375347 29474
rect 365732 29416 375286 29472
rect 375342 29416 375347 29472
rect 365732 29414 375347 29416
rect 365732 29412 365738 29414
rect 375281 29411 375347 29414
rect 386321 29338 386387 29341
rect 583520 29338 584960 29428
rect 386321 29336 393330 29338
rect 386321 29280 386326 29336
rect 386382 29280 393330 29336
rect 386321 29278 393330 29280
rect 386321 29275 386387 29278
rect 341566 29142 346410 29202
rect 360285 29202 360351 29205
rect 365662 29202 365668 29204
rect 360285 29200 365668 29202
rect 360285 29144 360290 29200
rect 360346 29144 365668 29200
rect 360285 29142 365668 29144
rect 360285 29139 360351 29142
rect 365662 29140 365668 29142
rect 365732 29140 365738 29204
rect 379421 29202 379487 29205
rect 376710 29200 379487 29202
rect 376710 29144 379426 29200
rect 379482 29144 379487 29200
rect 376710 29142 379487 29144
rect 393270 29202 393330 29278
rect 403022 29278 412650 29338
rect 393270 29142 402898 29202
rect 254485 29064 322122 29066
rect 254485 29008 254490 29064
rect 254546 29008 322122 29064
rect 254485 29006 322122 29008
rect 355961 29066 356027 29069
rect 360101 29066 360167 29069
rect 355961 29064 360167 29066
rect 355961 29008 355966 29064
rect 356022 29008 360106 29064
rect 360162 29008 360167 29064
rect 355961 29006 360167 29008
rect 254485 29003 254551 29006
rect 355961 29003 356027 29006
rect 360101 29003 360167 29006
rect 375281 29066 375347 29069
rect 376710 29066 376770 29142
rect 379421 29139 379487 29142
rect 375281 29064 376770 29066
rect 375281 29008 375286 29064
rect 375342 29008 376770 29064
rect 375281 29006 376770 29008
rect 402838 29066 402898 29142
rect 403022 29066 403082 29278
rect 412590 29202 412650 29278
rect 422342 29278 431970 29338
rect 412590 29142 422218 29202
rect 402838 29006 403082 29066
rect 422158 29066 422218 29142
rect 422342 29066 422402 29278
rect 431910 29202 431970 29278
rect 441662 29278 451290 29338
rect 431910 29142 441538 29202
rect 422158 29006 422402 29066
rect 441478 29066 441538 29142
rect 441662 29066 441722 29278
rect 451230 29202 451290 29278
rect 460982 29278 470610 29338
rect 451230 29142 460858 29202
rect 441478 29006 441722 29066
rect 460798 29066 460858 29142
rect 460982 29066 461042 29278
rect 470550 29202 470610 29278
rect 480302 29278 489930 29338
rect 470550 29142 480178 29202
rect 460798 29006 461042 29066
rect 480118 29066 480178 29142
rect 480302 29066 480362 29278
rect 489870 29202 489930 29278
rect 499622 29278 509250 29338
rect 489870 29142 499498 29202
rect 480118 29006 480362 29066
rect 499438 29066 499498 29142
rect 499622 29066 499682 29278
rect 509190 29202 509250 29278
rect 518942 29278 528570 29338
rect 509190 29142 518818 29202
rect 499438 29006 499682 29066
rect 518758 29066 518818 29142
rect 518942 29066 519002 29278
rect 528510 29202 528570 29278
rect 538262 29278 547890 29338
rect 528510 29142 538138 29202
rect 518758 29006 519002 29066
rect 538078 29066 538138 29142
rect 538262 29066 538322 29278
rect 547830 29202 547890 29278
rect 557582 29278 567210 29338
rect 547830 29142 557458 29202
rect 538078 29006 538322 29066
rect 557398 29066 557458 29142
rect 557582 29066 557642 29278
rect 567150 29202 567210 29278
rect 583342 29278 584960 29338
rect 583342 29202 583402 29278
rect 567150 29142 576778 29202
rect 557398 29006 557642 29066
rect 576718 29066 576778 29142
rect 576902 29142 583402 29202
rect 583520 29188 584960 29278
rect 576902 29066 576962 29142
rect 576718 29006 576962 29066
rect 375281 29003 375347 29006
rect 253105 26210 253171 26213
rect 253289 26210 253355 26213
rect 253105 26208 253355 26210
rect 253105 26152 253110 26208
rect 253166 26152 253294 26208
rect 253350 26152 253355 26208
rect 253105 26150 253355 26152
rect 253105 26147 253171 26150
rect 253289 26147 253355 26150
rect -960 21450 480 21540
rect 2865 21450 2931 21453
rect -960 21448 2931 21450
rect -960 21392 2870 21448
rect 2926 21392 2931 21448
rect -960 21390 2931 21392
rect -960 21300 480 21390
rect 2865 21387 2931 21390
rect 282361 19274 282427 19277
rect 286685 19274 286751 19277
rect 282318 19272 282427 19274
rect 282318 19216 282366 19272
rect 282422 19216 282427 19272
rect 282318 19211 282427 19216
rect 286550 19272 286751 19274
rect 286550 19216 286690 19272
rect 286746 19216 286751 19272
rect 286550 19214 286751 19216
rect 282318 19138 282378 19211
rect 283557 19138 283623 19141
rect 282318 19136 283623 19138
rect 282318 19080 283562 19136
rect 283618 19080 283623 19136
rect 282318 19078 283623 19080
rect 286550 19138 286610 19214
rect 286685 19211 286751 19214
rect 288433 19138 288499 19141
rect 286550 19136 288499 19138
rect 286550 19080 288438 19136
rect 288494 19080 288499 19136
rect 286550 19078 288499 19080
rect 283557 19075 283623 19078
rect 288433 19075 288499 19078
rect 324446 17988 324452 18052
rect 324516 18050 324522 18052
rect 328821 18050 328887 18053
rect 324516 18048 328887 18050
rect 324516 17992 328826 18048
rect 328882 17992 328887 18048
rect 324516 17990 328887 17992
rect 324516 17988 324522 17990
rect 328821 17987 328887 17990
rect 305913 17778 305979 17781
rect 492673 17778 492739 17781
rect 305913 17776 492739 17778
rect 305913 17720 305918 17776
rect 305974 17720 492678 17776
rect 492734 17720 492739 17776
rect 305913 17718 492739 17720
rect 305913 17715 305979 17718
rect 492673 17715 492739 17718
rect 314193 17642 314259 17645
rect 534073 17642 534139 17645
rect 583520 17642 584960 17732
rect 314193 17640 534139 17642
rect 314193 17584 314198 17640
rect 314254 17584 534078 17640
rect 534134 17584 534139 17640
rect 314193 17582 534139 17584
rect 314193 17579 314259 17582
rect 534073 17579 534139 17582
rect 583342 17582 584960 17642
rect 315573 17506 315639 17509
rect 536833 17506 536899 17509
rect 315573 17504 536899 17506
rect 315573 17448 315578 17504
rect 315634 17448 536838 17504
rect 536894 17448 536899 17504
rect 315573 17446 536899 17448
rect 315573 17443 315639 17446
rect 536833 17443 536899 17446
rect 315481 17370 315547 17373
rect 540973 17370 541039 17373
rect 315481 17368 541039 17370
rect 315481 17312 315486 17368
rect 315542 17312 540978 17368
rect 541034 17312 541039 17368
rect 315481 17310 541039 17312
rect 315481 17307 315547 17310
rect 540973 17307 541039 17310
rect 71681 17234 71747 17237
rect 338389 17234 338455 17237
rect 71681 17232 338455 17234
rect 71681 17176 71686 17232
rect 71742 17176 338394 17232
rect 338450 17176 338455 17232
rect 71681 17174 338455 17176
rect 71681 17171 71747 17174
rect 338389 17171 338455 17174
rect 259453 17098 259519 17101
rect 268694 17098 268700 17100
rect 259453 17096 268700 17098
rect 259453 17040 259458 17096
rect 259514 17040 268700 17096
rect 259453 17038 268700 17040
rect 259453 17035 259519 17038
rect 268694 17036 268700 17038
rect 268764 17036 268770 17100
rect 292573 17098 292639 17101
rect 300853 17098 300919 17101
rect 495341 17098 495407 17101
rect 292573 17096 300919 17098
rect 292573 17040 292578 17096
rect 292634 17040 300858 17096
rect 300914 17040 300919 17096
rect 292573 17038 300919 17040
rect 292573 17035 292639 17038
rect 300853 17035 300919 17038
rect 492676 17096 495407 17098
rect 492676 17040 495346 17096
rect 495402 17040 495407 17096
rect 492676 17038 495407 17040
rect 300853 16962 300919 16965
rect 332501 16962 332567 16965
rect 333881 16962 333947 16965
rect 244966 16902 249810 16962
rect 229093 16826 229159 16829
rect 244966 16826 245026 16902
rect 229093 16824 245026 16826
rect 229093 16768 229098 16824
rect 229154 16768 245026 16824
rect 229093 16766 245026 16768
rect 249750 16826 249810 16902
rect 300853 16960 310346 16962
rect 300853 16904 300858 16960
rect 300914 16904 310346 16960
rect 300853 16902 310346 16904
rect 300853 16899 300919 16902
rect 292573 16826 292639 16829
rect 249750 16766 249994 16826
rect 229093 16763 229159 16766
rect 249934 16690 249994 16766
rect 274590 16766 287714 16826
rect 259453 16690 259519 16693
rect 249934 16688 259519 16690
rect 249934 16632 259458 16688
rect 259514 16632 259519 16688
rect 249934 16630 259519 16632
rect 259453 16627 259519 16630
rect 268878 16628 268884 16692
rect 268948 16690 268954 16692
rect 274590 16690 274650 16766
rect 268948 16630 274650 16690
rect 287654 16690 287714 16766
rect 292438 16824 292639 16826
rect 292438 16768 292578 16824
rect 292634 16768 292639 16824
rect 292438 16766 292639 16768
rect 292438 16690 292498 16766
rect 292573 16763 292639 16766
rect 287654 16630 292498 16690
rect 310286 16690 310346 16902
rect 332501 16960 333947 16962
rect 332501 16904 332506 16960
rect 332562 16904 333886 16960
rect 333942 16904 333947 16960
rect 332501 16902 333947 16904
rect 332501 16899 332567 16902
rect 333881 16899 333947 16902
rect 311985 16826 312051 16829
rect 322933 16826 322999 16829
rect 369761 16826 369827 16829
rect 311985 16824 322999 16826
rect 311985 16768 311990 16824
rect 312046 16768 322938 16824
rect 322994 16768 322999 16824
rect 311985 16766 322999 16768
rect 311985 16763 312051 16766
rect 322933 16763 322999 16766
rect 346350 16824 369827 16826
rect 346350 16768 369766 16824
rect 369822 16768 369827 16824
rect 346350 16766 369827 16768
rect 311893 16690 311959 16693
rect 310286 16688 311959 16690
rect 310286 16632 311898 16688
rect 311954 16632 311959 16688
rect 310286 16630 311959 16632
rect 268948 16628 268954 16630
rect 311893 16627 311959 16630
rect 333881 16690 333947 16693
rect 336958 16690 336964 16692
rect 333881 16688 336964 16690
rect 333881 16632 333886 16688
rect 333942 16632 336964 16688
rect 333881 16630 336964 16632
rect 333881 16627 333947 16630
rect 336958 16628 336964 16630
rect 337028 16628 337034 16692
rect 346350 16557 346410 16766
rect 369761 16763 369827 16766
rect 379605 16826 379671 16829
rect 389081 16826 389147 16829
rect 379605 16824 389147 16826
rect 379605 16768 379610 16824
rect 379666 16768 389086 16824
rect 389142 16768 389147 16824
rect 379605 16766 389147 16768
rect 379605 16763 379671 16766
rect 389081 16763 389147 16766
rect 404261 16826 404327 16829
rect 408401 16826 408467 16829
rect 447041 16826 447107 16829
rect 404261 16824 408467 16826
rect 404261 16768 404266 16824
rect 404322 16768 408406 16824
rect 408462 16768 408467 16824
rect 404261 16766 408467 16768
rect 404261 16763 404327 16766
rect 408401 16763 408467 16766
rect 414016 16766 433442 16826
rect 369945 16690 370011 16693
rect 379421 16690 379487 16693
rect 369945 16688 379487 16690
rect 369945 16632 369950 16688
rect 370006 16632 379426 16688
rect 379482 16632 379487 16688
rect 369945 16630 379487 16632
rect 369945 16627 370011 16630
rect 379421 16627 379487 16630
rect 389265 16690 389331 16693
rect 394693 16690 394759 16693
rect 389265 16688 394759 16690
rect 389265 16632 389270 16688
rect 389326 16632 394698 16688
rect 394754 16632 394759 16688
rect 389265 16630 394759 16632
rect 389265 16627 389331 16630
rect 394693 16627 394759 16630
rect 408585 16690 408651 16693
rect 414016 16690 414076 16766
rect 408585 16688 414076 16690
rect 408585 16632 408590 16688
rect 408646 16632 414076 16688
rect 408585 16630 414076 16632
rect 433382 16690 433442 16766
rect 442950 16824 447107 16826
rect 442950 16768 447046 16824
rect 447102 16768 447107 16824
rect 442950 16766 447107 16768
rect 442950 16693 443010 16766
rect 447041 16763 447107 16766
rect 447225 16826 447291 16829
rect 466361 16826 466427 16829
rect 447225 16824 466427 16826
rect 447225 16768 447230 16824
rect 447286 16768 466366 16824
rect 466422 16768 466427 16824
rect 447225 16766 466427 16768
rect 447225 16763 447291 16766
rect 466361 16763 466427 16766
rect 476205 16826 476271 16829
rect 481582 16826 481588 16828
rect 476205 16824 481588 16826
rect 476205 16768 476210 16824
rect 476266 16768 481588 16824
rect 476205 16766 481588 16768
rect 476205 16763 476271 16766
rect 481582 16764 481588 16766
rect 481652 16764 481658 16828
rect 491201 16826 491267 16829
rect 492676 16826 492736 17038
rect 495341 17035 495407 17038
rect 495525 17098 495591 17101
rect 502374 17098 502380 17100
rect 495525 17096 502380 17098
rect 495525 17040 495530 17096
rect 495586 17040 502380 17096
rect 495525 17038 502380 17040
rect 495525 17035 495591 17038
rect 502374 17036 502380 17038
rect 502444 17036 502450 17100
rect 502374 16900 502380 16964
rect 502444 16962 502450 16964
rect 505001 16962 505067 16965
rect 502444 16960 505067 16962
rect 502444 16904 505006 16960
rect 505062 16904 505067 16960
rect 502444 16902 505067 16904
rect 502444 16900 502450 16902
rect 505001 16899 505067 16902
rect 518942 16902 528570 16962
rect 491201 16824 492736 16826
rect 491201 16768 491206 16824
rect 491262 16768 492736 16824
rect 491201 16766 492736 16768
rect 511901 16826 511967 16829
rect 511901 16824 518818 16826
rect 511901 16768 511906 16824
rect 511962 16768 518818 16824
rect 511901 16766 518818 16768
rect 491201 16763 491267 16766
rect 511901 16763 511967 16766
rect 437381 16690 437447 16693
rect 442901 16690 443010 16693
rect 433382 16688 437447 16690
rect 433382 16632 437386 16688
rect 437442 16632 437447 16688
rect 433382 16630 437447 16632
rect 442820 16688 443010 16690
rect 442820 16632 442906 16688
rect 442962 16632 443010 16688
rect 442820 16630 443010 16632
rect 466545 16690 466611 16693
rect 476021 16690 476087 16693
rect 466545 16688 476087 16690
rect 466545 16632 466550 16688
rect 466606 16632 476026 16688
rect 476082 16632 476087 16688
rect 466545 16630 476087 16632
rect 518758 16690 518818 16766
rect 518942 16690 519002 16902
rect 528510 16826 528570 16902
rect 538262 16902 547890 16962
rect 528510 16766 538138 16826
rect 518758 16630 519002 16690
rect 538078 16690 538138 16766
rect 538262 16690 538322 16902
rect 547830 16826 547890 16902
rect 557582 16902 567210 16962
rect 547830 16766 557458 16826
rect 538078 16630 538322 16690
rect 557398 16690 557458 16766
rect 557582 16690 557642 16902
rect 567150 16826 567210 16902
rect 583342 16826 583402 17582
rect 583520 17492 584960 17582
rect 567150 16766 576778 16826
rect 557398 16630 557642 16690
rect 576718 16690 576778 16766
rect 576902 16766 583402 16826
rect 576902 16690 576962 16766
rect 576718 16630 576962 16690
rect 408585 16627 408651 16630
rect 437381 16627 437447 16630
rect 442901 16627 442967 16630
rect 466545 16627 466611 16630
rect 476021 16627 476087 16630
rect 27521 16554 27587 16557
rect 278497 16554 278563 16557
rect 27521 16552 278563 16554
rect 27521 16496 27526 16552
rect 27582 16496 278502 16552
rect 278558 16496 278563 16552
rect 27521 16494 278563 16496
rect 27521 16491 27587 16494
rect 278497 16491 278563 16494
rect 278681 16554 278747 16557
rect 324262 16554 324268 16556
rect 278681 16552 324268 16554
rect 278681 16496 278686 16552
rect 278742 16496 324268 16552
rect 278681 16494 324268 16496
rect 278681 16491 278747 16494
rect 324262 16492 324268 16494
rect 324332 16492 324338 16556
rect 346350 16552 346459 16557
rect 346350 16496 346398 16552
rect 346454 16496 346459 16552
rect 346350 16494 346459 16496
rect 346393 16491 346459 16494
rect 481582 16492 481588 16556
rect 481652 16554 481658 16556
rect 491201 16554 491267 16557
rect 481652 16552 491267 16554
rect 481652 16496 491206 16552
rect 491262 16496 491267 16552
rect 481652 16494 491267 16496
rect 481652 16492 481658 16494
rect 491201 16491 491267 16494
rect 21909 16418 21975 16421
rect 268653 16418 268719 16421
rect 21909 16416 268719 16418
rect 21909 16360 21914 16416
rect 21970 16360 268658 16416
rect 268714 16360 268719 16416
rect 21909 16358 268719 16360
rect 21909 16355 21975 16358
rect 268653 16355 268719 16358
rect 269021 16418 269087 16421
rect 327349 16418 327415 16421
rect 269021 16416 327415 16418
rect 269021 16360 269026 16416
rect 269082 16360 327354 16416
rect 327410 16360 327415 16416
rect 269021 16358 327415 16360
rect 269021 16355 269087 16358
rect 327349 16355 327415 16358
rect 17861 16282 17927 16285
rect 264237 16282 264303 16285
rect 17861 16280 264303 16282
rect 17861 16224 17866 16280
rect 17922 16224 264242 16280
rect 264298 16224 264303 16280
rect 17861 16222 264303 16224
rect 17861 16219 17927 16222
rect 264237 16219 264303 16222
rect 268878 16220 268884 16284
rect 268948 16282 268954 16284
rect 278129 16282 278195 16285
rect 268948 16280 278195 16282
rect 268948 16224 278134 16280
rect 278190 16224 278195 16280
rect 268948 16222 278195 16224
rect 268948 16220 268954 16222
rect 278129 16219 278195 16222
rect 278681 16282 278747 16285
rect 297357 16282 297423 16285
rect 278681 16280 297423 16282
rect 278681 16224 278686 16280
rect 278742 16224 297362 16280
rect 297418 16224 297423 16280
rect 278681 16222 297423 16224
rect 278681 16219 278747 16222
rect 297357 16219 297423 16222
rect 301998 16220 302004 16284
rect 302068 16282 302074 16284
rect 308397 16282 308463 16285
rect 302068 16280 308463 16282
rect 302068 16224 308402 16280
rect 308458 16224 308463 16280
rect 302068 16222 308463 16224
rect 302068 16220 302074 16222
rect 308397 16219 308463 16222
rect 313038 16220 313044 16284
rect 313108 16282 313114 16284
rect 327441 16282 327507 16285
rect 313108 16280 327507 16282
rect 313108 16224 327446 16280
rect 327502 16224 327507 16280
rect 313108 16222 327507 16224
rect 313108 16220 313114 16222
rect 327441 16219 327507 16222
rect 336958 16220 336964 16284
rect 337028 16282 337034 16284
rect 345013 16282 345079 16285
rect 337028 16280 345079 16282
rect 337028 16224 345018 16280
rect 345074 16224 345079 16280
rect 337028 16222 345079 16224
rect 337028 16220 337034 16222
rect 345013 16219 345079 16222
rect 13721 16146 13787 16149
rect 325877 16146 325943 16149
rect 13721 16144 325943 16146
rect 13721 16088 13726 16144
rect 13782 16088 325882 16144
rect 325938 16088 325943 16144
rect 13721 16086 325943 16088
rect 13721 16083 13787 16086
rect 325877 16083 325943 16086
rect 9581 16010 9647 16013
rect 326153 16010 326219 16013
rect 9581 16008 326219 16010
rect 9581 15952 9586 16008
rect 9642 15952 326158 16008
rect 326214 15952 326219 16008
rect 9581 15950 326219 15952
rect 9581 15947 9647 15950
rect 326153 15947 326219 15950
rect 4061 15874 4127 15877
rect 324589 15874 324655 15877
rect 4061 15872 324655 15874
rect 4061 15816 4066 15872
rect 4122 15816 324594 15872
rect 324650 15816 324655 15872
rect 4061 15814 324655 15816
rect 4061 15811 4127 15814
rect 324589 15811 324655 15814
rect 264237 15602 264303 15605
rect 268878 15602 268884 15604
rect 264237 15600 268884 15602
rect 264237 15544 264242 15600
rect 264298 15544 268884 15600
rect 264237 15542 268884 15544
rect 264237 15539 264303 15542
rect 268878 15540 268884 15542
rect 268948 15540 268954 15604
rect 297357 15602 297423 15605
rect 301998 15602 302004 15604
rect 297357 15600 302004 15602
rect 297357 15544 297362 15600
rect 297418 15544 302004 15600
rect 297357 15542 302004 15544
rect 297357 15539 297423 15542
rect 301998 15540 302004 15542
rect 302068 15540 302074 15604
rect 308397 15602 308463 15605
rect 313038 15602 313044 15604
rect 308397 15600 313044 15602
rect 308397 15544 308402 15600
rect 308458 15544 313044 15600
rect 308397 15542 313044 15544
rect 308397 15539 308463 15542
rect 313038 15540 313044 15542
rect 313108 15540 313114 15604
rect 59261 15194 59327 15197
rect 335629 15194 335695 15197
rect 59261 15192 335695 15194
rect 59261 15136 59266 15192
rect 59322 15136 335634 15192
rect 335690 15136 335695 15192
rect 59261 15134 335695 15136
rect 59261 15131 59327 15134
rect 335629 15131 335695 15134
rect 56409 15058 56475 15061
rect 334525 15058 334591 15061
rect 56409 15056 334591 15058
rect 56409 15000 56414 15056
rect 56470 15000 334530 15056
rect 334586 15000 334591 15056
rect 56409 14998 334591 15000
rect 56409 14995 56475 14998
rect 334525 14995 334591 14998
rect 52361 14922 52427 14925
rect 334157 14922 334223 14925
rect 52361 14920 334223 14922
rect 52361 14864 52366 14920
rect 52422 14864 334162 14920
rect 334218 14864 334223 14920
rect 52361 14862 334223 14864
rect 52361 14859 52427 14862
rect 334157 14859 334223 14862
rect 48221 14786 48287 14789
rect 333237 14786 333303 14789
rect 48221 14784 333303 14786
rect 48221 14728 48226 14784
rect 48282 14728 333242 14784
rect 333298 14728 333303 14784
rect 48221 14726 333303 14728
rect 48221 14723 48287 14726
rect 333237 14723 333303 14726
rect 13629 14650 13695 14653
rect 325785 14650 325851 14653
rect 13629 14648 325851 14650
rect 13629 14592 13634 14648
rect 13690 14592 325790 14648
rect 325846 14592 325851 14648
rect 13629 14590 325851 14592
rect 13629 14587 13695 14590
rect 325785 14587 325851 14590
rect 8201 14514 8267 14517
rect 324773 14514 324839 14517
rect 8201 14512 324839 14514
rect 8201 14456 8206 14512
rect 8262 14456 324778 14512
rect 324834 14456 324839 14512
rect 8201 14454 324839 14456
rect 8201 14451 8267 14454
rect 324773 14451 324839 14454
rect 289353 13698 289419 13701
rect 414013 13698 414079 13701
rect 289353 13696 414079 13698
rect 289353 13640 289358 13696
rect 289414 13640 414018 13696
rect 414074 13640 414079 13696
rect 289353 13638 414079 13640
rect 289353 13635 289419 13638
rect 414013 13635 414079 13638
rect 290641 13562 290707 13565
rect 416773 13562 416839 13565
rect 290641 13560 416839 13562
rect 290641 13504 290646 13560
rect 290702 13504 416778 13560
rect 416834 13504 416839 13560
rect 290641 13502 416839 13504
rect 290641 13499 290707 13502
rect 416773 13499 416839 13502
rect 290825 13426 290891 13429
rect 420913 13426 420979 13429
rect 290825 13424 420979 13426
rect 290825 13368 290830 13424
rect 290886 13368 420918 13424
rect 420974 13368 420979 13424
rect 290825 13366 420979 13368
rect 290825 13363 290891 13366
rect 420913 13363 420979 13366
rect 291929 13290 291995 13293
rect 425053 13290 425119 13293
rect 291929 13288 425119 13290
rect 291929 13232 291934 13288
rect 291990 13232 425058 13288
rect 425114 13232 425119 13288
rect 291929 13230 425119 13232
rect 291929 13227 291995 13230
rect 425053 13227 425119 13230
rect 292113 13154 292179 13157
rect 427813 13154 427879 13157
rect 292113 13152 427879 13154
rect 292113 13096 292118 13152
rect 292174 13096 427818 13152
rect 427874 13096 427879 13152
rect 292113 13094 427879 13096
rect 292113 13091 292179 13094
rect 427813 13091 427879 13094
rect 3969 13018 4035 13021
rect 324405 13018 324471 13021
rect 3969 13016 324471 13018
rect 3969 12960 3974 13016
rect 4030 12960 324410 13016
rect 324466 12960 324471 13016
rect 3969 12958 324471 12960
rect 3969 12955 4035 12958
rect 324405 12955 324471 12958
rect 319713 12338 319779 12341
rect 560293 12338 560359 12341
rect 319713 12336 560359 12338
rect 319713 12280 319718 12336
rect 319774 12280 560298 12336
rect 560354 12280 560359 12336
rect 319713 12278 560359 12280
rect 319713 12275 319779 12278
rect 560293 12275 560359 12278
rect 319529 12202 319595 12205
rect 563053 12202 563119 12205
rect 319529 12200 563119 12202
rect 319529 12144 319534 12200
rect 319590 12144 563058 12200
rect 563114 12144 563119 12200
rect 319529 12142 563119 12144
rect 319529 12139 319595 12142
rect 563053 12139 563119 12142
rect 321001 12066 321067 12069
rect 567193 12066 567259 12069
rect 321001 12064 567259 12066
rect 321001 12008 321006 12064
rect 321062 12008 567198 12064
rect 567254 12008 567259 12064
rect 321001 12006 567259 12008
rect 321001 12003 321067 12006
rect 567193 12003 567259 12006
rect 322289 11930 322355 11933
rect 574093 11930 574159 11933
rect 322289 11928 574159 11930
rect 322289 11872 322294 11928
rect 322350 11872 574098 11928
rect 574154 11872 574159 11928
rect 322289 11870 574159 11872
rect 322289 11867 322355 11870
rect 574093 11867 574159 11870
rect 2681 11794 2747 11797
rect 323301 11794 323367 11797
rect 2681 11792 323367 11794
rect 2681 11736 2686 11792
rect 2742 11736 323306 11792
rect 323362 11736 323367 11792
rect 2681 11734 323367 11736
rect 2681 11731 2747 11734
rect 323301 11731 323367 11734
rect 323945 11794 324011 11797
rect 578233 11794 578299 11797
rect 323945 11792 578299 11794
rect 323945 11736 323950 11792
rect 324006 11736 578238 11792
rect 578294 11736 578299 11792
rect 323945 11734 578299 11736
rect 323945 11731 324011 11734
rect 578233 11731 578299 11734
rect 1301 11658 1367 11661
rect 323393 11658 323459 11661
rect 1301 11656 323459 11658
rect 1301 11600 1306 11656
rect 1362 11600 323398 11656
rect 323454 11600 323459 11656
rect 1301 11598 323459 11600
rect 1301 11595 1367 11598
rect 323393 11595 323459 11598
rect 324037 11658 324103 11661
rect 580993 11658 581059 11661
rect 324037 11656 581059 11658
rect 324037 11600 324042 11656
rect 324098 11600 580998 11656
rect 581054 11600 581059 11656
rect 324037 11598 581059 11600
rect 324037 11595 324103 11598
rect 580993 11595 581059 11598
rect 322473 11250 322539 11253
rect 322430 11248 322539 11250
rect 322430 11192 322478 11248
rect 322534 11192 322539 11248
rect 322430 11187 322539 11192
rect 322430 10978 322490 11187
rect 328637 10978 328703 10981
rect 322430 10976 328703 10978
rect 322430 10920 328642 10976
rect 328698 10920 328703 10976
rect 322430 10918 328703 10920
rect 328637 10915 328703 10918
rect 300485 10842 300551 10845
rect 466453 10842 466519 10845
rect 300485 10840 466519 10842
rect 300485 10784 300490 10840
rect 300546 10784 466458 10840
rect 466514 10784 466519 10840
rect 300485 10782 466519 10784
rect 300485 10779 300551 10782
rect 466453 10779 466519 10782
rect 300577 10706 300643 10709
rect 469213 10706 469279 10709
rect 300577 10704 469279 10706
rect 300577 10648 300582 10704
rect 300638 10648 469218 10704
rect 469274 10648 469279 10704
rect 300577 10646 469279 10648
rect 300577 10643 300643 10646
rect 469213 10643 469279 10646
rect 301957 10570 302023 10573
rect 473353 10570 473419 10573
rect 301957 10568 473419 10570
rect 301957 10512 301962 10568
rect 302018 10512 473358 10568
rect 473414 10512 473419 10568
rect 301957 10510 473419 10512
rect 301957 10507 302023 10510
rect 473353 10507 473419 10510
rect 303429 10434 303495 10437
rect 477585 10434 477651 10437
rect 303429 10432 477651 10434
rect 303429 10376 303434 10432
rect 303490 10376 477590 10432
rect 477646 10376 477651 10432
rect 303429 10374 477651 10376
rect 303429 10371 303495 10374
rect 477585 10371 477651 10374
rect 303337 10298 303403 10301
rect 480253 10298 480319 10301
rect 303337 10296 480319 10298
rect 303337 10240 303342 10296
rect 303398 10240 480258 10296
rect 480314 10240 480319 10296
rect 303337 10238 480319 10240
rect 303337 10235 303403 10238
rect 480253 10235 480319 10238
rect 100477 9754 100543 9757
rect 100661 9754 100727 9757
rect 100477 9752 100727 9754
rect 100477 9696 100482 9752
rect 100538 9696 100666 9752
rect 100722 9696 100727 9752
rect 100477 9694 100727 9696
rect 100477 9691 100543 9694
rect 100661 9691 100727 9694
rect 284109 9618 284175 9621
rect 384665 9618 384731 9621
rect 284109 9616 384731 9618
rect 284109 9560 284114 9616
rect 284170 9560 384670 9616
rect 384726 9560 384731 9616
rect 284109 9558 384731 9560
rect 284109 9555 284175 9558
rect 384665 9555 384731 9558
rect 317137 9482 317203 9485
rect 548885 9482 548951 9485
rect 317137 9480 548951 9482
rect 317137 9424 317142 9480
rect 317198 9424 548890 9480
rect 548946 9424 548951 9480
rect 317137 9422 548951 9424
rect 317137 9419 317203 9422
rect 548885 9419 548951 9422
rect 318425 9346 318491 9349
rect 555969 9346 556035 9349
rect 318425 9344 556035 9346
rect 318425 9288 318430 9344
rect 318486 9288 555974 9344
rect 556030 9288 556035 9344
rect 318425 9286 556035 9288
rect 318425 9283 318491 9286
rect 555969 9283 556035 9286
rect 319805 9210 319871 9213
rect 559557 9210 559623 9213
rect 319805 9208 559623 9210
rect 319805 9152 319810 9208
rect 319866 9152 559562 9208
rect 559618 9152 559623 9208
rect 319805 9150 559623 9152
rect 319805 9147 319871 9150
rect 559557 9147 559623 9150
rect 319897 9074 319963 9077
rect 563145 9074 563211 9077
rect 319897 9072 563211 9074
rect 319897 9016 319902 9072
rect 319958 9016 563150 9072
rect 563206 9016 563211 9072
rect 319897 9014 563211 9016
rect 319897 9011 319963 9014
rect 563145 9011 563211 9014
rect 321185 8938 321251 8941
rect 570229 8938 570295 8941
rect 321185 8936 570295 8938
rect 321185 8880 321190 8936
rect 321246 8880 570234 8936
rect 570290 8880 570295 8936
rect 321185 8878 570295 8880
rect 321185 8875 321251 8878
rect 570229 8875 570295 8878
rect 150433 8258 150499 8261
rect 234889 8258 234955 8261
rect 150433 8256 234955 8258
rect 150433 8200 150438 8256
rect 150494 8200 234894 8256
rect 234950 8200 234955 8256
rect 150433 8198 234955 8200
rect 150433 8195 150499 8198
rect 234889 8195 234955 8198
rect 308765 8258 308831 8261
rect 509601 8258 509667 8261
rect 308765 8256 509667 8258
rect 308765 8200 308770 8256
rect 308826 8200 509606 8256
rect 509662 8200 509667 8256
rect 308765 8198 509667 8200
rect 308765 8195 308831 8198
rect 509601 8195 509667 8198
rect 146845 8122 146911 8125
rect 233509 8122 233575 8125
rect 146845 8120 233575 8122
rect 146845 8064 146850 8120
rect 146906 8064 233514 8120
rect 233570 8064 233575 8120
rect 146845 8062 233575 8064
rect 146845 8059 146911 8062
rect 233509 8059 233575 8062
rect 310237 8122 310303 8125
rect 513189 8122 513255 8125
rect 310237 8120 513255 8122
rect 310237 8064 310242 8120
rect 310298 8064 513194 8120
rect 513250 8064 513255 8120
rect 310237 8062 513255 8064
rect 310237 8059 310303 8062
rect 513189 8059 513255 8062
rect 143257 7986 143323 7989
rect 233417 7986 233483 7989
rect 143257 7984 233483 7986
rect 143257 7928 143262 7984
rect 143318 7928 233422 7984
rect 233478 7928 233483 7984
rect 143257 7926 233483 7928
rect 143257 7923 143323 7926
rect 233417 7923 233483 7926
rect 310145 7986 310211 7989
rect 516777 7986 516843 7989
rect 310145 7984 516843 7986
rect 310145 7928 310150 7984
rect 310206 7928 516782 7984
rect 516838 7928 516843 7984
rect 310145 7926 516843 7928
rect 310145 7923 310211 7926
rect 516777 7923 516843 7926
rect 139669 7850 139735 7853
rect 232313 7850 232379 7853
rect 139669 7848 232379 7850
rect 139669 7792 139674 7848
rect 139730 7792 232318 7848
rect 232374 7792 232379 7848
rect 139669 7790 232379 7792
rect 139669 7787 139735 7790
rect 232313 7787 232379 7790
rect 311525 7850 311591 7853
rect 523861 7850 523927 7853
rect 311525 7848 523927 7850
rect 311525 7792 311530 7848
rect 311586 7792 523866 7848
rect 523922 7792 523927 7848
rect 311525 7790 523927 7792
rect 311525 7787 311591 7790
rect 523861 7787 523927 7790
rect 136081 7714 136147 7717
rect 232221 7714 232287 7717
rect 136081 7712 232287 7714
rect 136081 7656 136086 7712
rect 136142 7656 232226 7712
rect 232282 7656 232287 7712
rect 136081 7654 232287 7656
rect 136081 7651 136147 7654
rect 232221 7651 232287 7654
rect 312905 7714 312971 7717
rect 527449 7714 527515 7717
rect 312905 7712 527515 7714
rect 312905 7656 312910 7712
rect 312966 7656 527454 7712
rect 527510 7656 527515 7712
rect 312905 7654 527515 7656
rect 312905 7651 312971 7654
rect 527449 7651 527515 7654
rect 132585 7578 132651 7581
rect 230841 7578 230907 7581
rect 132585 7576 230907 7578
rect 132585 7520 132590 7576
rect 132646 7520 230846 7576
rect 230902 7520 230907 7576
rect 132585 7518 230907 7520
rect 132585 7515 132651 7518
rect 230841 7515 230907 7518
rect 312997 7578 313063 7581
rect 531037 7578 531103 7581
rect 312997 7576 531103 7578
rect 312997 7520 313002 7576
rect 313058 7520 531042 7576
rect 531098 7520 531103 7576
rect 312997 7518 531103 7520
rect 312997 7515 313063 7518
rect 531037 7515 531103 7518
rect -960 7170 480 7260
rect 3417 7170 3483 7173
rect -960 7168 3483 7170
rect -960 7112 3422 7168
rect 3478 7112 3483 7168
rect -960 7110 3483 7112
rect -960 7020 480 7110
rect 3417 7107 3483 7110
rect 149237 6898 149303 6901
rect 234797 6898 234863 6901
rect 149237 6896 234863 6898
rect 149237 6840 149242 6896
rect 149298 6840 234802 6896
rect 234858 6840 234863 6896
rect 149237 6838 234863 6840
rect 149237 6835 149303 6838
rect 234797 6835 234863 6838
rect 321277 6898 321343 6901
rect 327073 6898 327139 6901
rect 321277 6896 327139 6898
rect 321277 6840 321282 6896
rect 321338 6840 327078 6896
rect 327134 6840 327139 6896
rect 321277 6838 327139 6840
rect 321277 6835 321343 6838
rect 327073 6835 327139 6838
rect 145649 6762 145715 6765
rect 233693 6762 233759 6765
rect 145649 6760 233759 6762
rect 145649 6704 145654 6760
rect 145710 6704 233698 6760
rect 233754 6704 233759 6760
rect 145649 6702 233759 6704
rect 145649 6699 145715 6702
rect 233693 6699 233759 6702
rect 289629 6762 289695 6765
rect 415669 6762 415735 6765
rect 289629 6760 415735 6762
rect 289629 6704 289634 6760
rect 289690 6704 415674 6760
rect 415730 6704 415735 6760
rect 289629 6702 415735 6704
rect 289629 6699 289695 6702
rect 415669 6699 415735 6702
rect 142061 6626 142127 6629
rect 232589 6626 232655 6629
rect 142061 6624 232655 6626
rect 142061 6568 142066 6624
rect 142122 6568 232594 6624
rect 232650 6568 232655 6624
rect 142061 6566 232655 6568
rect 142061 6563 142127 6566
rect 232589 6563 232655 6566
rect 291009 6626 291075 6629
rect 419165 6626 419231 6629
rect 291009 6624 419231 6626
rect 291009 6568 291014 6624
rect 291070 6568 419170 6624
rect 419226 6568 419231 6624
rect 291009 6566 419231 6568
rect 291009 6563 291075 6566
rect 419165 6563 419231 6566
rect 138473 6490 138539 6493
rect 232037 6490 232103 6493
rect 138473 6488 232103 6490
rect 138473 6432 138478 6488
rect 138534 6432 232042 6488
rect 232098 6432 232103 6488
rect 138473 6430 232103 6432
rect 138473 6427 138539 6430
rect 232037 6427 232103 6430
rect 291101 6490 291167 6493
rect 422753 6490 422819 6493
rect 291101 6488 422819 6490
rect 291101 6432 291106 6488
rect 291162 6432 422758 6488
rect 422814 6432 422819 6488
rect 291101 6430 422819 6432
rect 291101 6427 291167 6430
rect 422753 6427 422819 6430
rect 134885 6354 134951 6357
rect 231209 6354 231275 6357
rect 134885 6352 231275 6354
rect 134885 6296 134890 6352
rect 134946 6296 231214 6352
rect 231270 6296 231275 6352
rect 134885 6294 231275 6296
rect 134885 6291 134951 6294
rect 231209 6291 231275 6294
rect 292389 6354 292455 6357
rect 426341 6354 426407 6357
rect 292389 6352 426407 6354
rect 292389 6296 292394 6352
rect 292450 6296 426346 6352
rect 426402 6296 426407 6352
rect 292389 6294 426407 6296
rect 292389 6291 292455 6294
rect 426341 6291 426407 6294
rect 131389 6218 131455 6221
rect 230749 6218 230815 6221
rect 131389 6216 230815 6218
rect 131389 6160 131394 6216
rect 131450 6160 230754 6216
rect 230810 6160 230815 6216
rect 131389 6158 230815 6160
rect 131389 6155 131455 6158
rect 230749 6155 230815 6158
rect 292481 6218 292547 6221
rect 429929 6218 429995 6221
rect 292481 6216 429995 6218
rect 292481 6160 292486 6216
rect 292542 6160 429934 6216
rect 429990 6160 429995 6216
rect 292481 6158 429995 6160
rect 292481 6155 292547 6158
rect 429929 6155 429995 6158
rect 583520 5796 584960 6036
rect 205081 5538 205147 5541
rect 245745 5538 245811 5541
rect 205081 5536 245811 5538
rect 205081 5480 205086 5536
rect 205142 5480 245750 5536
rect 245806 5480 245811 5536
rect 205081 5478 245811 5480
rect 205081 5475 205147 5478
rect 245745 5475 245811 5478
rect 267549 5538 267615 5541
rect 309777 5538 309843 5541
rect 267549 5536 309843 5538
rect 267549 5480 267554 5536
rect 267610 5480 309782 5536
rect 309838 5480 309843 5536
rect 267549 5478 309843 5480
rect 267549 5475 267615 5478
rect 309777 5475 309843 5478
rect 319989 5538 320055 5541
rect 561949 5538 562015 5541
rect 319989 5536 562015 5538
rect 319989 5480 319994 5536
rect 320050 5480 561954 5536
rect 562010 5480 562015 5536
rect 319989 5478 562015 5480
rect 319989 5475 320055 5478
rect 561949 5475 562015 5478
rect 190821 5402 190887 5405
rect 242893 5402 242959 5405
rect 190821 5400 242959 5402
rect 190821 5344 190826 5400
rect 190882 5344 242898 5400
rect 242954 5344 242959 5400
rect 190821 5342 242959 5344
rect 190821 5339 190887 5342
rect 242893 5339 242959 5342
rect 269021 5402 269087 5405
rect 313365 5402 313431 5405
rect 269021 5400 313431 5402
rect 269021 5344 269026 5400
rect 269082 5344 313370 5400
rect 313426 5344 313431 5400
rect 269021 5342 313431 5344
rect 269021 5339 269087 5342
rect 313365 5339 313431 5342
rect 321369 5402 321435 5405
rect 565537 5402 565603 5405
rect 321369 5400 565603 5402
rect 321369 5344 321374 5400
rect 321430 5344 565542 5400
rect 565598 5344 565603 5400
rect 321369 5342 565603 5344
rect 321369 5339 321435 5342
rect 565537 5339 565603 5342
rect 183737 5266 183803 5269
rect 242065 5266 242131 5269
rect 183737 5264 242131 5266
rect 183737 5208 183742 5264
rect 183798 5208 242070 5264
rect 242126 5208 242131 5264
rect 183737 5206 242131 5208
rect 183737 5203 183803 5206
rect 242065 5203 242131 5206
rect 270217 5266 270283 5269
rect 317045 5266 317111 5269
rect 270217 5264 317111 5266
rect 270217 5208 270222 5264
rect 270278 5208 317050 5264
rect 317106 5208 317111 5264
rect 270217 5206 317111 5208
rect 270217 5203 270283 5206
rect 317045 5203 317111 5206
rect 321461 5266 321527 5269
rect 569033 5266 569099 5269
rect 321461 5264 569099 5266
rect 321461 5208 321466 5264
rect 321522 5208 569038 5264
rect 569094 5208 569099 5264
rect 321461 5206 569099 5208
rect 321461 5203 321527 5206
rect 569033 5203 569099 5206
rect 176561 5130 176627 5133
rect 240133 5130 240199 5133
rect 176561 5128 240199 5130
rect 176561 5072 176566 5128
rect 176622 5072 240138 5128
rect 240194 5072 240199 5128
rect 176561 5070 240199 5072
rect 176561 5067 176627 5070
rect 240133 5067 240199 5070
rect 268837 5130 268903 5133
rect 315757 5130 315823 5133
rect 268837 5128 315823 5130
rect 268837 5072 268842 5128
rect 268898 5072 315762 5128
rect 315818 5072 315823 5128
rect 268837 5070 315823 5072
rect 268837 5067 268903 5070
rect 315757 5067 315823 5070
rect 322657 5130 322723 5133
rect 572621 5130 572687 5133
rect 322657 5128 572687 5130
rect 322657 5072 322662 5128
rect 322718 5072 572626 5128
rect 572682 5072 572687 5128
rect 322657 5070 572687 5072
rect 322657 5067 322723 5070
rect 572621 5067 572687 5070
rect 137277 4994 137343 4997
rect 231853 4994 231919 4997
rect 137277 4992 231919 4994
rect 137277 4936 137282 4992
rect 137338 4936 231858 4992
rect 231914 4936 231919 4992
rect 137277 4934 231919 4936
rect 137277 4931 137343 4934
rect 231853 4931 231919 4934
rect 270401 4994 270467 4997
rect 319253 4994 319319 4997
rect 270401 4992 319319 4994
rect 270401 4936 270406 4992
rect 270462 4936 319258 4992
rect 319314 4936 319319 4992
rect 270401 4934 319319 4936
rect 270401 4931 270467 4934
rect 319253 4931 319319 4934
rect 322841 4994 322907 4997
rect 576209 4994 576275 4997
rect 322841 4992 576275 4994
rect 322841 4936 322846 4992
rect 322902 4936 576214 4992
rect 576270 4936 576275 4992
rect 322841 4934 576275 4936
rect 322841 4931 322907 4934
rect 576209 4931 576275 4934
rect 130193 4858 130259 4861
rect 230565 4858 230631 4861
rect 130193 4856 230631 4858
rect 130193 4800 130198 4856
rect 130254 4800 230570 4856
rect 230626 4800 230631 4856
rect 130193 4798 230631 4800
rect 130193 4795 130259 4798
rect 230565 4795 230631 4798
rect 270309 4858 270375 4861
rect 322841 4858 322907 4861
rect 270309 4856 322907 4858
rect 270309 4800 270314 4856
rect 270370 4800 322846 4856
rect 322902 4800 322907 4856
rect 270309 4798 322907 4800
rect 270309 4795 270375 4798
rect 322841 4795 322907 4798
rect 324221 4858 324287 4861
rect 579797 4858 579863 4861
rect 324221 4856 579863 4858
rect 324221 4800 324226 4856
rect 324282 4800 579802 4856
rect 579858 4800 579863 4856
rect 324221 4798 579863 4800
rect 324221 4795 324287 4798
rect 579797 4795 579863 4798
rect 273069 4178 273135 4181
rect 273345 4178 273411 4181
rect 273069 4176 273411 4178
rect 273069 4120 273074 4176
rect 273130 4120 273350 4176
rect 273406 4120 273411 4176
rect 273069 4118 273411 4120
rect 273069 4115 273135 4118
rect 273345 4115 273411 4118
rect 292389 4178 292455 4181
rect 292665 4178 292731 4181
rect 292389 4176 292731 4178
rect 292389 4120 292394 4176
rect 292450 4120 292670 4176
rect 292726 4120 292731 4176
rect 292389 4118 292731 4120
rect 292389 4115 292455 4118
rect 292665 4115 292731 4118
rect 311801 4178 311867 4181
rect 313917 4178 313983 4181
rect 311801 4176 313983 4178
rect 311801 4120 311806 4176
rect 311862 4120 313922 4176
rect 313978 4120 313983 4176
rect 311801 4118 313983 4120
rect 311801 4115 311867 4118
rect 313917 4115 313983 4118
rect 324865 4178 324931 4181
rect 330293 4178 330359 4181
rect 324865 4176 330359 4178
rect 324865 4120 324870 4176
rect 324926 4120 330298 4176
rect 330354 4120 330359 4176
rect 324865 4118 330359 4120
rect 324865 4115 324931 4118
rect 330293 4115 330359 4118
rect 24301 4042 24367 4045
rect 328545 4042 328611 4045
rect 24301 4040 328611 4042
rect 24301 3984 24306 4040
rect 24362 3984 328550 4040
rect 328606 3984 328611 4040
rect 24301 3982 328611 3984
rect 24301 3979 24367 3982
rect 328545 3979 328611 3982
rect 23105 3906 23171 3909
rect 328729 3906 328795 3909
rect 23105 3904 328795 3906
rect 23105 3848 23110 3904
rect 23166 3848 328734 3904
rect 328790 3848 328795 3904
rect 23105 3846 328795 3848
rect 23105 3843 23171 3846
rect 328729 3843 328795 3846
rect 18321 3770 18387 3773
rect 327257 3770 327323 3773
rect 18321 3768 327323 3770
rect 18321 3712 18326 3768
rect 18382 3712 327262 3768
rect 327318 3712 327323 3768
rect 18321 3710 327323 3712
rect 18321 3707 18387 3710
rect 327257 3707 327323 3710
rect 16021 3634 16087 3637
rect 327533 3634 327599 3637
rect 16021 3632 327599 3634
rect 16021 3576 16026 3632
rect 16082 3576 327538 3632
rect 327594 3576 327599 3632
rect 16021 3574 327599 3576
rect 16021 3571 16087 3574
rect 327533 3571 327599 3574
rect 14825 3498 14891 3501
rect 326061 3498 326127 3501
rect 14825 3496 326127 3498
rect 14825 3440 14830 3496
rect 14886 3440 326066 3496
rect 326122 3440 326127 3496
rect 14825 3438 326127 3440
rect 14825 3435 14891 3438
rect 326061 3435 326127 3438
rect 6453 3362 6519 3365
rect 324313 3362 324379 3365
rect 6453 3360 324379 3362
rect 6453 3304 6458 3360
rect 6514 3304 324318 3360
rect 324374 3304 324379 3360
rect 6453 3302 324379 3304
rect 6453 3299 6519 3302
rect 324313 3299 324379 3302
rect 224769 3226 224835 3229
rect 224953 3226 225019 3229
rect 224769 3224 225019 3226
rect 224769 3168 224774 3224
rect 224830 3168 224958 3224
rect 225014 3168 225019 3224
rect 224769 3166 225019 3168
rect 224769 3163 224835 3166
rect 224953 3163 225019 3166
rect 263409 3226 263475 3229
rect 263685 3226 263751 3229
rect 263409 3224 263751 3226
rect 263409 3168 263414 3224
rect 263470 3168 263690 3224
rect 263746 3168 263751 3224
rect 263409 3166 263751 3168
rect 263409 3163 263475 3166
rect 263685 3163 263751 3166
rect 275185 3226 275251 3229
rect 282821 3226 282887 3229
rect 275185 3224 282887 3226
rect 275185 3168 275190 3224
rect 275246 3168 282826 3224
rect 282882 3168 282887 3224
rect 275185 3166 282887 3168
rect 275185 3163 275251 3166
rect 282821 3163 282887 3166
<< via3 >>
rect 348372 462980 348436 463044
rect 232452 462844 232516 462908
rect 348740 462708 348804 462772
rect 348924 462572 348988 462636
rect 348556 462436 348620 462500
rect 344324 459988 344388 460052
rect 344140 459852 344204 459916
rect 342484 459716 342548 459780
rect 231716 459640 231780 459644
rect 231716 459584 231730 459640
rect 231730 459584 231780 459640
rect 231716 459580 231780 459584
rect 233004 459580 233068 459644
rect 233924 459580 233988 459644
rect 342668 459580 342732 459644
rect 343588 459580 343652 459644
rect 345428 459580 345492 459644
rect 233740 459308 233804 459372
rect 258948 459308 259012 459372
rect 324636 459308 324700 459372
rect 345244 459308 345308 459372
rect 347084 459308 347148 459372
rect 258948 457812 259012 457876
rect 324636 457676 324700 457740
rect 232452 452508 232516 452572
rect 348924 415652 348988 415716
rect 348740 392260 348804 392324
rect 348556 368732 348620 368796
rect 348372 345340 348436 345404
rect 266492 337996 266556 338060
rect 266492 328476 266556 328540
rect 344324 310660 344388 310724
rect 376708 310796 376772 310860
rect 357388 310524 357452 310588
rect 376708 310524 376772 310588
rect 357388 310252 357452 310316
rect 344140 263740 344204 263804
rect 376708 263876 376772 263940
rect 357388 263604 357452 263668
rect 376708 263604 376772 263668
rect 357388 263332 357452 263396
rect 232084 220824 232148 220828
rect 232084 220768 232098 220824
rect 232098 220768 232148 220824
rect 232084 220764 232148 220768
rect 342484 216820 342548 216884
rect 376708 216956 376772 217020
rect 357388 216684 357452 216748
rect 376708 216684 376772 216748
rect 357388 216412 357452 216476
rect 232084 211168 232148 211172
rect 232084 211112 232098 211168
rect 232098 211112 232148 211168
rect 232084 211108 232148 211112
rect 342668 169900 342732 169964
rect 376708 170036 376772 170100
rect 357388 169764 357452 169828
rect 376708 169764 376772 169828
rect 357388 169492 357452 169556
rect 244412 138680 244476 138684
rect 244412 138624 244462 138680
rect 244462 138624 244476 138680
rect 244412 138620 244476 138624
rect 244412 125624 244476 125628
rect 244412 125568 244426 125624
rect 244426 125568 244476 125624
rect 244412 125564 244476 125568
rect 233740 90476 233804 90540
rect 365668 87348 365732 87412
rect 365668 87076 365732 87140
rect 343588 80004 343652 80068
rect 345244 64772 345308 64836
rect 324268 63956 324332 64020
rect 343588 63956 343652 64020
rect 233924 63684 233988 63748
rect 258028 63684 258092 63748
rect 315988 63684 316052 63748
rect 324268 63684 324332 63748
rect 343588 63684 343652 63748
rect 376708 63820 376772 63884
rect 258028 63412 258092 63476
rect 277164 63548 277228 63612
rect 376708 63548 376772 63612
rect 315988 63276 316052 63340
rect 277164 63140 277228 63204
rect 345428 50900 345492 50964
rect 237420 40428 237484 40492
rect 277164 40428 277228 40492
rect 277164 40020 277228 40084
rect 376708 40292 376772 40356
rect 231716 39884 231780 39948
rect 237420 39884 237484 39948
rect 357388 40020 357452 40084
rect 376708 40020 376772 40084
rect 357388 39748 357452 39812
rect 347084 35804 347148 35868
rect 241468 29412 241532 29476
rect 233004 29140 233068 29204
rect 241468 29140 241532 29204
rect 365668 29412 365732 29476
rect 365668 29140 365732 29204
rect 324452 17988 324516 18052
rect 268700 17036 268764 17100
rect 268884 16628 268948 16692
rect 336964 16628 337028 16692
rect 481588 16764 481652 16828
rect 502380 17036 502444 17100
rect 502380 16900 502444 16964
rect 324268 16492 324332 16556
rect 481588 16492 481652 16556
rect 268884 16220 268948 16284
rect 302004 16220 302068 16284
rect 313044 16220 313108 16284
rect 336964 16220 337028 16284
rect 268884 15540 268948 15604
rect 302004 15540 302068 15604
rect 313044 15540 313108 15604
<< metal4 >>
rect -8436 711278 -7836 711300
rect -8436 711042 -8254 711278
rect -8018 711042 -7836 711278
rect -8436 710958 -7836 711042
rect -8436 710722 -8254 710958
rect -8018 710722 -7836 710958
rect -8436 679254 -7836 710722
rect -8436 679018 -8254 679254
rect -8018 679018 -7836 679254
rect -8436 678934 -7836 679018
rect -8436 678698 -8254 678934
rect -8018 678698 -7836 678934
rect -8436 643254 -7836 678698
rect -8436 643018 -8254 643254
rect -8018 643018 -7836 643254
rect -8436 642934 -7836 643018
rect -8436 642698 -8254 642934
rect -8018 642698 -7836 642934
rect -8436 607254 -7836 642698
rect -8436 607018 -8254 607254
rect -8018 607018 -7836 607254
rect -8436 606934 -7836 607018
rect -8436 606698 -8254 606934
rect -8018 606698 -7836 606934
rect -8436 571254 -7836 606698
rect -8436 571018 -8254 571254
rect -8018 571018 -7836 571254
rect -8436 570934 -7836 571018
rect -8436 570698 -8254 570934
rect -8018 570698 -7836 570934
rect -8436 535254 -7836 570698
rect -8436 535018 -8254 535254
rect -8018 535018 -7836 535254
rect -8436 534934 -7836 535018
rect -8436 534698 -8254 534934
rect -8018 534698 -7836 534934
rect -8436 499254 -7836 534698
rect -8436 499018 -8254 499254
rect -8018 499018 -7836 499254
rect -8436 498934 -7836 499018
rect -8436 498698 -8254 498934
rect -8018 498698 -7836 498934
rect -8436 463254 -7836 498698
rect -8436 463018 -8254 463254
rect -8018 463018 -7836 463254
rect -8436 462934 -7836 463018
rect -8436 462698 -8254 462934
rect -8018 462698 -7836 462934
rect -8436 427254 -7836 462698
rect -8436 427018 -8254 427254
rect -8018 427018 -7836 427254
rect -8436 426934 -7836 427018
rect -8436 426698 -8254 426934
rect -8018 426698 -7836 426934
rect -8436 391254 -7836 426698
rect -8436 391018 -8254 391254
rect -8018 391018 -7836 391254
rect -8436 390934 -7836 391018
rect -8436 390698 -8254 390934
rect -8018 390698 -7836 390934
rect -8436 355254 -7836 390698
rect -8436 355018 -8254 355254
rect -8018 355018 -7836 355254
rect -8436 354934 -7836 355018
rect -8436 354698 -8254 354934
rect -8018 354698 -7836 354934
rect -8436 319254 -7836 354698
rect -8436 319018 -8254 319254
rect -8018 319018 -7836 319254
rect -8436 318934 -7836 319018
rect -8436 318698 -8254 318934
rect -8018 318698 -7836 318934
rect -8436 283254 -7836 318698
rect -8436 283018 -8254 283254
rect -8018 283018 -7836 283254
rect -8436 282934 -7836 283018
rect -8436 282698 -8254 282934
rect -8018 282698 -7836 282934
rect -8436 247254 -7836 282698
rect -8436 247018 -8254 247254
rect -8018 247018 -7836 247254
rect -8436 246934 -7836 247018
rect -8436 246698 -8254 246934
rect -8018 246698 -7836 246934
rect -8436 211254 -7836 246698
rect -8436 211018 -8254 211254
rect -8018 211018 -7836 211254
rect -8436 210934 -7836 211018
rect -8436 210698 -8254 210934
rect -8018 210698 -7836 210934
rect -8436 175254 -7836 210698
rect -8436 175018 -8254 175254
rect -8018 175018 -7836 175254
rect -8436 174934 -7836 175018
rect -8436 174698 -8254 174934
rect -8018 174698 -7836 174934
rect -8436 139254 -7836 174698
rect -8436 139018 -8254 139254
rect -8018 139018 -7836 139254
rect -8436 138934 -7836 139018
rect -8436 138698 -8254 138934
rect -8018 138698 -7836 138934
rect -8436 103254 -7836 138698
rect -8436 103018 -8254 103254
rect -8018 103018 -7836 103254
rect -8436 102934 -7836 103018
rect -8436 102698 -8254 102934
rect -8018 102698 -7836 102934
rect -8436 67254 -7836 102698
rect -8436 67018 -8254 67254
rect -8018 67018 -7836 67254
rect -8436 66934 -7836 67018
rect -8436 66698 -8254 66934
rect -8018 66698 -7836 66934
rect -8436 31254 -7836 66698
rect -8436 31018 -8254 31254
rect -8018 31018 -7836 31254
rect -8436 30934 -7836 31018
rect -8436 30698 -8254 30934
rect -8018 30698 -7836 30934
rect -8436 -6786 -7836 30698
rect -7516 710358 -6916 710380
rect -7516 710122 -7334 710358
rect -7098 710122 -6916 710358
rect -7516 710038 -6916 710122
rect -7516 709802 -7334 710038
rect -7098 709802 -6916 710038
rect -7516 697254 -6916 709802
rect 11604 710358 12204 711300
rect 11604 710122 11786 710358
rect 12022 710122 12204 710358
rect 11604 710038 12204 710122
rect 11604 709802 11786 710038
rect 12022 709802 12204 710038
rect -7516 697018 -7334 697254
rect -7098 697018 -6916 697254
rect -7516 696934 -6916 697018
rect -7516 696698 -7334 696934
rect -7098 696698 -6916 696934
rect -7516 661254 -6916 696698
rect -7516 661018 -7334 661254
rect -7098 661018 -6916 661254
rect -7516 660934 -6916 661018
rect -7516 660698 -7334 660934
rect -7098 660698 -6916 660934
rect -7516 625254 -6916 660698
rect -7516 625018 -7334 625254
rect -7098 625018 -6916 625254
rect -7516 624934 -6916 625018
rect -7516 624698 -7334 624934
rect -7098 624698 -6916 624934
rect -7516 589254 -6916 624698
rect -7516 589018 -7334 589254
rect -7098 589018 -6916 589254
rect -7516 588934 -6916 589018
rect -7516 588698 -7334 588934
rect -7098 588698 -6916 588934
rect -7516 553254 -6916 588698
rect -7516 553018 -7334 553254
rect -7098 553018 -6916 553254
rect -7516 552934 -6916 553018
rect -7516 552698 -7334 552934
rect -7098 552698 -6916 552934
rect -7516 517254 -6916 552698
rect -7516 517018 -7334 517254
rect -7098 517018 -6916 517254
rect -7516 516934 -6916 517018
rect -7516 516698 -7334 516934
rect -7098 516698 -6916 516934
rect -7516 481254 -6916 516698
rect -7516 481018 -7334 481254
rect -7098 481018 -6916 481254
rect -7516 480934 -6916 481018
rect -7516 480698 -7334 480934
rect -7098 480698 -6916 480934
rect -7516 445254 -6916 480698
rect -7516 445018 -7334 445254
rect -7098 445018 -6916 445254
rect -7516 444934 -6916 445018
rect -7516 444698 -7334 444934
rect -7098 444698 -6916 444934
rect -7516 409254 -6916 444698
rect -7516 409018 -7334 409254
rect -7098 409018 -6916 409254
rect -7516 408934 -6916 409018
rect -7516 408698 -7334 408934
rect -7098 408698 -6916 408934
rect -7516 373254 -6916 408698
rect -7516 373018 -7334 373254
rect -7098 373018 -6916 373254
rect -7516 372934 -6916 373018
rect -7516 372698 -7334 372934
rect -7098 372698 -6916 372934
rect -7516 337254 -6916 372698
rect -7516 337018 -7334 337254
rect -7098 337018 -6916 337254
rect -7516 336934 -6916 337018
rect -7516 336698 -7334 336934
rect -7098 336698 -6916 336934
rect -7516 301254 -6916 336698
rect -7516 301018 -7334 301254
rect -7098 301018 -6916 301254
rect -7516 300934 -6916 301018
rect -7516 300698 -7334 300934
rect -7098 300698 -6916 300934
rect -7516 265254 -6916 300698
rect -7516 265018 -7334 265254
rect -7098 265018 -6916 265254
rect -7516 264934 -6916 265018
rect -7516 264698 -7334 264934
rect -7098 264698 -6916 264934
rect -7516 229254 -6916 264698
rect -7516 229018 -7334 229254
rect -7098 229018 -6916 229254
rect -7516 228934 -6916 229018
rect -7516 228698 -7334 228934
rect -7098 228698 -6916 228934
rect -7516 193254 -6916 228698
rect -7516 193018 -7334 193254
rect -7098 193018 -6916 193254
rect -7516 192934 -6916 193018
rect -7516 192698 -7334 192934
rect -7098 192698 -6916 192934
rect -7516 157254 -6916 192698
rect -7516 157018 -7334 157254
rect -7098 157018 -6916 157254
rect -7516 156934 -6916 157018
rect -7516 156698 -7334 156934
rect -7098 156698 -6916 156934
rect -7516 121254 -6916 156698
rect -7516 121018 -7334 121254
rect -7098 121018 -6916 121254
rect -7516 120934 -6916 121018
rect -7516 120698 -7334 120934
rect -7098 120698 -6916 120934
rect -7516 85254 -6916 120698
rect -7516 85018 -7334 85254
rect -7098 85018 -6916 85254
rect -7516 84934 -6916 85018
rect -7516 84698 -7334 84934
rect -7098 84698 -6916 84934
rect -7516 49254 -6916 84698
rect -7516 49018 -7334 49254
rect -7098 49018 -6916 49254
rect -7516 48934 -6916 49018
rect -7516 48698 -7334 48934
rect -7098 48698 -6916 48934
rect -7516 13254 -6916 48698
rect -7516 13018 -7334 13254
rect -7098 13018 -6916 13254
rect -7516 12934 -6916 13018
rect -7516 12698 -7334 12934
rect -7098 12698 -6916 12934
rect -7516 -5866 -6916 12698
rect -6596 709438 -5996 709460
rect -6596 709202 -6414 709438
rect -6178 709202 -5996 709438
rect -6596 709118 -5996 709202
rect -6596 708882 -6414 709118
rect -6178 708882 -5996 709118
rect -6596 675654 -5996 708882
rect -6596 675418 -6414 675654
rect -6178 675418 -5996 675654
rect -6596 675334 -5996 675418
rect -6596 675098 -6414 675334
rect -6178 675098 -5996 675334
rect -6596 639654 -5996 675098
rect -6596 639418 -6414 639654
rect -6178 639418 -5996 639654
rect -6596 639334 -5996 639418
rect -6596 639098 -6414 639334
rect -6178 639098 -5996 639334
rect -6596 603654 -5996 639098
rect -6596 603418 -6414 603654
rect -6178 603418 -5996 603654
rect -6596 603334 -5996 603418
rect -6596 603098 -6414 603334
rect -6178 603098 -5996 603334
rect -6596 567654 -5996 603098
rect -6596 567418 -6414 567654
rect -6178 567418 -5996 567654
rect -6596 567334 -5996 567418
rect -6596 567098 -6414 567334
rect -6178 567098 -5996 567334
rect -6596 531654 -5996 567098
rect -6596 531418 -6414 531654
rect -6178 531418 -5996 531654
rect -6596 531334 -5996 531418
rect -6596 531098 -6414 531334
rect -6178 531098 -5996 531334
rect -6596 495654 -5996 531098
rect -6596 495418 -6414 495654
rect -6178 495418 -5996 495654
rect -6596 495334 -5996 495418
rect -6596 495098 -6414 495334
rect -6178 495098 -5996 495334
rect -6596 459654 -5996 495098
rect -6596 459418 -6414 459654
rect -6178 459418 -5996 459654
rect -6596 459334 -5996 459418
rect -6596 459098 -6414 459334
rect -6178 459098 -5996 459334
rect -6596 423654 -5996 459098
rect -6596 423418 -6414 423654
rect -6178 423418 -5996 423654
rect -6596 423334 -5996 423418
rect -6596 423098 -6414 423334
rect -6178 423098 -5996 423334
rect -6596 387654 -5996 423098
rect -6596 387418 -6414 387654
rect -6178 387418 -5996 387654
rect -6596 387334 -5996 387418
rect -6596 387098 -6414 387334
rect -6178 387098 -5996 387334
rect -6596 351654 -5996 387098
rect -6596 351418 -6414 351654
rect -6178 351418 -5996 351654
rect -6596 351334 -5996 351418
rect -6596 351098 -6414 351334
rect -6178 351098 -5996 351334
rect -6596 315654 -5996 351098
rect -6596 315418 -6414 315654
rect -6178 315418 -5996 315654
rect -6596 315334 -5996 315418
rect -6596 315098 -6414 315334
rect -6178 315098 -5996 315334
rect -6596 279654 -5996 315098
rect -6596 279418 -6414 279654
rect -6178 279418 -5996 279654
rect -6596 279334 -5996 279418
rect -6596 279098 -6414 279334
rect -6178 279098 -5996 279334
rect -6596 243654 -5996 279098
rect -6596 243418 -6414 243654
rect -6178 243418 -5996 243654
rect -6596 243334 -5996 243418
rect -6596 243098 -6414 243334
rect -6178 243098 -5996 243334
rect -6596 207654 -5996 243098
rect -6596 207418 -6414 207654
rect -6178 207418 -5996 207654
rect -6596 207334 -5996 207418
rect -6596 207098 -6414 207334
rect -6178 207098 -5996 207334
rect -6596 171654 -5996 207098
rect -6596 171418 -6414 171654
rect -6178 171418 -5996 171654
rect -6596 171334 -5996 171418
rect -6596 171098 -6414 171334
rect -6178 171098 -5996 171334
rect -6596 135654 -5996 171098
rect -6596 135418 -6414 135654
rect -6178 135418 -5996 135654
rect -6596 135334 -5996 135418
rect -6596 135098 -6414 135334
rect -6178 135098 -5996 135334
rect -6596 99654 -5996 135098
rect -6596 99418 -6414 99654
rect -6178 99418 -5996 99654
rect -6596 99334 -5996 99418
rect -6596 99098 -6414 99334
rect -6178 99098 -5996 99334
rect -6596 63654 -5996 99098
rect -6596 63418 -6414 63654
rect -6178 63418 -5996 63654
rect -6596 63334 -5996 63418
rect -6596 63098 -6414 63334
rect -6178 63098 -5996 63334
rect -6596 27654 -5996 63098
rect -6596 27418 -6414 27654
rect -6178 27418 -5996 27654
rect -6596 27334 -5996 27418
rect -6596 27098 -6414 27334
rect -6178 27098 -5996 27334
rect -6596 -4946 -5996 27098
rect -5676 708518 -5076 708540
rect -5676 708282 -5494 708518
rect -5258 708282 -5076 708518
rect -5676 708198 -5076 708282
rect -5676 707962 -5494 708198
rect -5258 707962 -5076 708198
rect -5676 693654 -5076 707962
rect 8004 708518 8604 709460
rect 8004 708282 8186 708518
rect 8422 708282 8604 708518
rect 8004 708198 8604 708282
rect 8004 707962 8186 708198
rect 8422 707962 8604 708198
rect -5676 693418 -5494 693654
rect -5258 693418 -5076 693654
rect -5676 693334 -5076 693418
rect -5676 693098 -5494 693334
rect -5258 693098 -5076 693334
rect -5676 657654 -5076 693098
rect -5676 657418 -5494 657654
rect -5258 657418 -5076 657654
rect -5676 657334 -5076 657418
rect -5676 657098 -5494 657334
rect -5258 657098 -5076 657334
rect -5676 621654 -5076 657098
rect -5676 621418 -5494 621654
rect -5258 621418 -5076 621654
rect -5676 621334 -5076 621418
rect -5676 621098 -5494 621334
rect -5258 621098 -5076 621334
rect -5676 585654 -5076 621098
rect -5676 585418 -5494 585654
rect -5258 585418 -5076 585654
rect -5676 585334 -5076 585418
rect -5676 585098 -5494 585334
rect -5258 585098 -5076 585334
rect -5676 549654 -5076 585098
rect -5676 549418 -5494 549654
rect -5258 549418 -5076 549654
rect -5676 549334 -5076 549418
rect -5676 549098 -5494 549334
rect -5258 549098 -5076 549334
rect -5676 513654 -5076 549098
rect -5676 513418 -5494 513654
rect -5258 513418 -5076 513654
rect -5676 513334 -5076 513418
rect -5676 513098 -5494 513334
rect -5258 513098 -5076 513334
rect -5676 477654 -5076 513098
rect -5676 477418 -5494 477654
rect -5258 477418 -5076 477654
rect -5676 477334 -5076 477418
rect -5676 477098 -5494 477334
rect -5258 477098 -5076 477334
rect -5676 441654 -5076 477098
rect -5676 441418 -5494 441654
rect -5258 441418 -5076 441654
rect -5676 441334 -5076 441418
rect -5676 441098 -5494 441334
rect -5258 441098 -5076 441334
rect -5676 405654 -5076 441098
rect -5676 405418 -5494 405654
rect -5258 405418 -5076 405654
rect -5676 405334 -5076 405418
rect -5676 405098 -5494 405334
rect -5258 405098 -5076 405334
rect -5676 369654 -5076 405098
rect -5676 369418 -5494 369654
rect -5258 369418 -5076 369654
rect -5676 369334 -5076 369418
rect -5676 369098 -5494 369334
rect -5258 369098 -5076 369334
rect -5676 333654 -5076 369098
rect -5676 333418 -5494 333654
rect -5258 333418 -5076 333654
rect -5676 333334 -5076 333418
rect -5676 333098 -5494 333334
rect -5258 333098 -5076 333334
rect -5676 297654 -5076 333098
rect -5676 297418 -5494 297654
rect -5258 297418 -5076 297654
rect -5676 297334 -5076 297418
rect -5676 297098 -5494 297334
rect -5258 297098 -5076 297334
rect -5676 261654 -5076 297098
rect -5676 261418 -5494 261654
rect -5258 261418 -5076 261654
rect -5676 261334 -5076 261418
rect -5676 261098 -5494 261334
rect -5258 261098 -5076 261334
rect -5676 225654 -5076 261098
rect -5676 225418 -5494 225654
rect -5258 225418 -5076 225654
rect -5676 225334 -5076 225418
rect -5676 225098 -5494 225334
rect -5258 225098 -5076 225334
rect -5676 189654 -5076 225098
rect -5676 189418 -5494 189654
rect -5258 189418 -5076 189654
rect -5676 189334 -5076 189418
rect -5676 189098 -5494 189334
rect -5258 189098 -5076 189334
rect -5676 153654 -5076 189098
rect -5676 153418 -5494 153654
rect -5258 153418 -5076 153654
rect -5676 153334 -5076 153418
rect -5676 153098 -5494 153334
rect -5258 153098 -5076 153334
rect -5676 117654 -5076 153098
rect -5676 117418 -5494 117654
rect -5258 117418 -5076 117654
rect -5676 117334 -5076 117418
rect -5676 117098 -5494 117334
rect -5258 117098 -5076 117334
rect -5676 81654 -5076 117098
rect -5676 81418 -5494 81654
rect -5258 81418 -5076 81654
rect -5676 81334 -5076 81418
rect -5676 81098 -5494 81334
rect -5258 81098 -5076 81334
rect -5676 45654 -5076 81098
rect -5676 45418 -5494 45654
rect -5258 45418 -5076 45654
rect -5676 45334 -5076 45418
rect -5676 45098 -5494 45334
rect -5258 45098 -5076 45334
rect -5676 9654 -5076 45098
rect -5676 9418 -5494 9654
rect -5258 9418 -5076 9654
rect -5676 9334 -5076 9418
rect -5676 9098 -5494 9334
rect -5258 9098 -5076 9334
rect -5676 -4026 -5076 9098
rect -4756 707598 -4156 707620
rect -4756 707362 -4574 707598
rect -4338 707362 -4156 707598
rect -4756 707278 -4156 707362
rect -4756 707042 -4574 707278
rect -4338 707042 -4156 707278
rect -4756 672054 -4156 707042
rect -4756 671818 -4574 672054
rect -4338 671818 -4156 672054
rect -4756 671734 -4156 671818
rect -4756 671498 -4574 671734
rect -4338 671498 -4156 671734
rect -4756 636054 -4156 671498
rect -4756 635818 -4574 636054
rect -4338 635818 -4156 636054
rect -4756 635734 -4156 635818
rect -4756 635498 -4574 635734
rect -4338 635498 -4156 635734
rect -4756 600054 -4156 635498
rect -4756 599818 -4574 600054
rect -4338 599818 -4156 600054
rect -4756 599734 -4156 599818
rect -4756 599498 -4574 599734
rect -4338 599498 -4156 599734
rect -4756 564054 -4156 599498
rect -4756 563818 -4574 564054
rect -4338 563818 -4156 564054
rect -4756 563734 -4156 563818
rect -4756 563498 -4574 563734
rect -4338 563498 -4156 563734
rect -4756 528054 -4156 563498
rect -4756 527818 -4574 528054
rect -4338 527818 -4156 528054
rect -4756 527734 -4156 527818
rect -4756 527498 -4574 527734
rect -4338 527498 -4156 527734
rect -4756 492054 -4156 527498
rect -4756 491818 -4574 492054
rect -4338 491818 -4156 492054
rect -4756 491734 -4156 491818
rect -4756 491498 -4574 491734
rect -4338 491498 -4156 491734
rect -4756 456054 -4156 491498
rect -4756 455818 -4574 456054
rect -4338 455818 -4156 456054
rect -4756 455734 -4156 455818
rect -4756 455498 -4574 455734
rect -4338 455498 -4156 455734
rect -4756 420054 -4156 455498
rect -4756 419818 -4574 420054
rect -4338 419818 -4156 420054
rect -4756 419734 -4156 419818
rect -4756 419498 -4574 419734
rect -4338 419498 -4156 419734
rect -4756 384054 -4156 419498
rect -4756 383818 -4574 384054
rect -4338 383818 -4156 384054
rect -4756 383734 -4156 383818
rect -4756 383498 -4574 383734
rect -4338 383498 -4156 383734
rect -4756 348054 -4156 383498
rect -4756 347818 -4574 348054
rect -4338 347818 -4156 348054
rect -4756 347734 -4156 347818
rect -4756 347498 -4574 347734
rect -4338 347498 -4156 347734
rect -4756 312054 -4156 347498
rect -4756 311818 -4574 312054
rect -4338 311818 -4156 312054
rect -4756 311734 -4156 311818
rect -4756 311498 -4574 311734
rect -4338 311498 -4156 311734
rect -4756 276054 -4156 311498
rect -4756 275818 -4574 276054
rect -4338 275818 -4156 276054
rect -4756 275734 -4156 275818
rect -4756 275498 -4574 275734
rect -4338 275498 -4156 275734
rect -4756 240054 -4156 275498
rect -4756 239818 -4574 240054
rect -4338 239818 -4156 240054
rect -4756 239734 -4156 239818
rect -4756 239498 -4574 239734
rect -4338 239498 -4156 239734
rect -4756 204054 -4156 239498
rect -4756 203818 -4574 204054
rect -4338 203818 -4156 204054
rect -4756 203734 -4156 203818
rect -4756 203498 -4574 203734
rect -4338 203498 -4156 203734
rect -4756 168054 -4156 203498
rect -4756 167818 -4574 168054
rect -4338 167818 -4156 168054
rect -4756 167734 -4156 167818
rect -4756 167498 -4574 167734
rect -4338 167498 -4156 167734
rect -4756 132054 -4156 167498
rect -4756 131818 -4574 132054
rect -4338 131818 -4156 132054
rect -4756 131734 -4156 131818
rect -4756 131498 -4574 131734
rect -4338 131498 -4156 131734
rect -4756 96054 -4156 131498
rect -4756 95818 -4574 96054
rect -4338 95818 -4156 96054
rect -4756 95734 -4156 95818
rect -4756 95498 -4574 95734
rect -4338 95498 -4156 95734
rect -4756 60054 -4156 95498
rect -4756 59818 -4574 60054
rect -4338 59818 -4156 60054
rect -4756 59734 -4156 59818
rect -4756 59498 -4574 59734
rect -4338 59498 -4156 59734
rect -4756 24054 -4156 59498
rect -4756 23818 -4574 24054
rect -4338 23818 -4156 24054
rect -4756 23734 -4156 23818
rect -4756 23498 -4574 23734
rect -4338 23498 -4156 23734
rect -4756 -3106 -4156 23498
rect -3836 706678 -3236 706700
rect -3836 706442 -3654 706678
rect -3418 706442 -3236 706678
rect -3836 706358 -3236 706442
rect -3836 706122 -3654 706358
rect -3418 706122 -3236 706358
rect -3836 690054 -3236 706122
rect 4404 706678 5004 707620
rect 4404 706442 4586 706678
rect 4822 706442 5004 706678
rect 4404 706358 5004 706442
rect 4404 706122 4586 706358
rect 4822 706122 5004 706358
rect -3836 689818 -3654 690054
rect -3418 689818 -3236 690054
rect -3836 689734 -3236 689818
rect -3836 689498 -3654 689734
rect -3418 689498 -3236 689734
rect -3836 654054 -3236 689498
rect -3836 653818 -3654 654054
rect -3418 653818 -3236 654054
rect -3836 653734 -3236 653818
rect -3836 653498 -3654 653734
rect -3418 653498 -3236 653734
rect -3836 618054 -3236 653498
rect -3836 617818 -3654 618054
rect -3418 617818 -3236 618054
rect -3836 617734 -3236 617818
rect -3836 617498 -3654 617734
rect -3418 617498 -3236 617734
rect -3836 582054 -3236 617498
rect -3836 581818 -3654 582054
rect -3418 581818 -3236 582054
rect -3836 581734 -3236 581818
rect -3836 581498 -3654 581734
rect -3418 581498 -3236 581734
rect -3836 546054 -3236 581498
rect -3836 545818 -3654 546054
rect -3418 545818 -3236 546054
rect -3836 545734 -3236 545818
rect -3836 545498 -3654 545734
rect -3418 545498 -3236 545734
rect -3836 510054 -3236 545498
rect -3836 509818 -3654 510054
rect -3418 509818 -3236 510054
rect -3836 509734 -3236 509818
rect -3836 509498 -3654 509734
rect -3418 509498 -3236 509734
rect -3836 474054 -3236 509498
rect -3836 473818 -3654 474054
rect -3418 473818 -3236 474054
rect -3836 473734 -3236 473818
rect -3836 473498 -3654 473734
rect -3418 473498 -3236 473734
rect -3836 438054 -3236 473498
rect -3836 437818 -3654 438054
rect -3418 437818 -3236 438054
rect -3836 437734 -3236 437818
rect -3836 437498 -3654 437734
rect -3418 437498 -3236 437734
rect -3836 402054 -3236 437498
rect -3836 401818 -3654 402054
rect -3418 401818 -3236 402054
rect -3836 401734 -3236 401818
rect -3836 401498 -3654 401734
rect -3418 401498 -3236 401734
rect -3836 366054 -3236 401498
rect -3836 365818 -3654 366054
rect -3418 365818 -3236 366054
rect -3836 365734 -3236 365818
rect -3836 365498 -3654 365734
rect -3418 365498 -3236 365734
rect -3836 330054 -3236 365498
rect -3836 329818 -3654 330054
rect -3418 329818 -3236 330054
rect -3836 329734 -3236 329818
rect -3836 329498 -3654 329734
rect -3418 329498 -3236 329734
rect -3836 294054 -3236 329498
rect -3836 293818 -3654 294054
rect -3418 293818 -3236 294054
rect -3836 293734 -3236 293818
rect -3836 293498 -3654 293734
rect -3418 293498 -3236 293734
rect -3836 258054 -3236 293498
rect -3836 257818 -3654 258054
rect -3418 257818 -3236 258054
rect -3836 257734 -3236 257818
rect -3836 257498 -3654 257734
rect -3418 257498 -3236 257734
rect -3836 222054 -3236 257498
rect -3836 221818 -3654 222054
rect -3418 221818 -3236 222054
rect -3836 221734 -3236 221818
rect -3836 221498 -3654 221734
rect -3418 221498 -3236 221734
rect -3836 186054 -3236 221498
rect -3836 185818 -3654 186054
rect -3418 185818 -3236 186054
rect -3836 185734 -3236 185818
rect -3836 185498 -3654 185734
rect -3418 185498 -3236 185734
rect -3836 150054 -3236 185498
rect -3836 149818 -3654 150054
rect -3418 149818 -3236 150054
rect -3836 149734 -3236 149818
rect -3836 149498 -3654 149734
rect -3418 149498 -3236 149734
rect -3836 114054 -3236 149498
rect -3836 113818 -3654 114054
rect -3418 113818 -3236 114054
rect -3836 113734 -3236 113818
rect -3836 113498 -3654 113734
rect -3418 113498 -3236 113734
rect -3836 78054 -3236 113498
rect -3836 77818 -3654 78054
rect -3418 77818 -3236 78054
rect -3836 77734 -3236 77818
rect -3836 77498 -3654 77734
rect -3418 77498 -3236 77734
rect -3836 42054 -3236 77498
rect -3836 41818 -3654 42054
rect -3418 41818 -3236 42054
rect -3836 41734 -3236 41818
rect -3836 41498 -3654 41734
rect -3418 41498 -3236 41734
rect -3836 6054 -3236 41498
rect -3836 5818 -3654 6054
rect -3418 5818 -3236 6054
rect -3836 5734 -3236 5818
rect -3836 5498 -3654 5734
rect -3418 5498 -3236 5734
rect -3836 -2186 -3236 5498
rect -2916 705758 -2316 705780
rect -2916 705522 -2734 705758
rect -2498 705522 -2316 705758
rect -2916 705438 -2316 705522
rect -2916 705202 -2734 705438
rect -2498 705202 -2316 705438
rect -2916 668454 -2316 705202
rect -2916 668218 -2734 668454
rect -2498 668218 -2316 668454
rect -2916 668134 -2316 668218
rect -2916 667898 -2734 668134
rect -2498 667898 -2316 668134
rect -2916 632454 -2316 667898
rect -2916 632218 -2734 632454
rect -2498 632218 -2316 632454
rect -2916 632134 -2316 632218
rect -2916 631898 -2734 632134
rect -2498 631898 -2316 632134
rect -2916 596454 -2316 631898
rect -2916 596218 -2734 596454
rect -2498 596218 -2316 596454
rect -2916 596134 -2316 596218
rect -2916 595898 -2734 596134
rect -2498 595898 -2316 596134
rect -2916 560454 -2316 595898
rect -2916 560218 -2734 560454
rect -2498 560218 -2316 560454
rect -2916 560134 -2316 560218
rect -2916 559898 -2734 560134
rect -2498 559898 -2316 560134
rect -2916 524454 -2316 559898
rect -2916 524218 -2734 524454
rect -2498 524218 -2316 524454
rect -2916 524134 -2316 524218
rect -2916 523898 -2734 524134
rect -2498 523898 -2316 524134
rect -2916 488454 -2316 523898
rect -2916 488218 -2734 488454
rect -2498 488218 -2316 488454
rect -2916 488134 -2316 488218
rect -2916 487898 -2734 488134
rect -2498 487898 -2316 488134
rect -2916 452454 -2316 487898
rect -2916 452218 -2734 452454
rect -2498 452218 -2316 452454
rect -2916 452134 -2316 452218
rect -2916 451898 -2734 452134
rect -2498 451898 -2316 452134
rect -2916 416454 -2316 451898
rect -2916 416218 -2734 416454
rect -2498 416218 -2316 416454
rect -2916 416134 -2316 416218
rect -2916 415898 -2734 416134
rect -2498 415898 -2316 416134
rect -2916 380454 -2316 415898
rect -2916 380218 -2734 380454
rect -2498 380218 -2316 380454
rect -2916 380134 -2316 380218
rect -2916 379898 -2734 380134
rect -2498 379898 -2316 380134
rect -2916 344454 -2316 379898
rect -2916 344218 -2734 344454
rect -2498 344218 -2316 344454
rect -2916 344134 -2316 344218
rect -2916 343898 -2734 344134
rect -2498 343898 -2316 344134
rect -2916 308454 -2316 343898
rect -2916 308218 -2734 308454
rect -2498 308218 -2316 308454
rect -2916 308134 -2316 308218
rect -2916 307898 -2734 308134
rect -2498 307898 -2316 308134
rect -2916 272454 -2316 307898
rect -2916 272218 -2734 272454
rect -2498 272218 -2316 272454
rect -2916 272134 -2316 272218
rect -2916 271898 -2734 272134
rect -2498 271898 -2316 272134
rect -2916 236454 -2316 271898
rect -2916 236218 -2734 236454
rect -2498 236218 -2316 236454
rect -2916 236134 -2316 236218
rect -2916 235898 -2734 236134
rect -2498 235898 -2316 236134
rect -2916 200454 -2316 235898
rect -2916 200218 -2734 200454
rect -2498 200218 -2316 200454
rect -2916 200134 -2316 200218
rect -2916 199898 -2734 200134
rect -2498 199898 -2316 200134
rect -2916 164454 -2316 199898
rect -2916 164218 -2734 164454
rect -2498 164218 -2316 164454
rect -2916 164134 -2316 164218
rect -2916 163898 -2734 164134
rect -2498 163898 -2316 164134
rect -2916 128454 -2316 163898
rect -2916 128218 -2734 128454
rect -2498 128218 -2316 128454
rect -2916 128134 -2316 128218
rect -2916 127898 -2734 128134
rect -2498 127898 -2316 128134
rect -2916 92454 -2316 127898
rect -2916 92218 -2734 92454
rect -2498 92218 -2316 92454
rect -2916 92134 -2316 92218
rect -2916 91898 -2734 92134
rect -2498 91898 -2316 92134
rect -2916 56454 -2316 91898
rect -2916 56218 -2734 56454
rect -2498 56218 -2316 56454
rect -2916 56134 -2316 56218
rect -2916 55898 -2734 56134
rect -2498 55898 -2316 56134
rect -2916 20454 -2316 55898
rect -2916 20218 -2734 20454
rect -2498 20218 -2316 20454
rect -2916 20134 -2316 20218
rect -2916 19898 -2734 20134
rect -2498 19898 -2316 20134
rect -2916 -1266 -2316 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705780
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2916 -1502 -2734 -1266
rect -2498 -1502 -2316 -1266
rect -2916 -1586 -2316 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 -2316 -1586
rect -2916 -1844 -2316 -1822
rect 804 -1844 1404 -902
rect 4404 690054 5004 706122
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3836 -2422 -3654 -2186
rect -3418 -2422 -3236 -2186
rect -3836 -2506 -3236 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 -3236 -2506
rect -3836 -2764 -3236 -2742
rect 4404 -2186 5004 5498
rect 4404 -2422 4586 -2186
rect 4822 -2422 5004 -2186
rect 4404 -2506 5004 -2422
rect 4404 -2742 4586 -2506
rect 4822 -2742 5004 -2506
rect -4756 -3342 -4574 -3106
rect -4338 -3342 -4156 -3106
rect -4756 -3426 -4156 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 -4156 -3426
rect -4756 -3684 -4156 -3662
rect 4404 -3684 5004 -2742
rect 8004 693654 8604 707962
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5676 -4262 -5494 -4026
rect -5258 -4262 -5076 -4026
rect -5676 -4346 -5076 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 -5076 -4346
rect -5676 -4604 -5076 -4582
rect 8004 -4026 8604 9098
rect 8004 -4262 8186 -4026
rect 8422 -4262 8604 -4026
rect 8004 -4346 8604 -4262
rect 8004 -4582 8186 -4346
rect 8422 -4582 8604 -4346
rect -6596 -5182 -6414 -4946
rect -6178 -5182 -5996 -4946
rect -6596 -5266 -5996 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 -5996 -5266
rect -6596 -5524 -5996 -5502
rect 8004 -5524 8604 -4582
rect 11604 697254 12204 709802
rect 29604 711278 30204 711300
rect 29604 711042 29786 711278
rect 30022 711042 30204 711278
rect 29604 710958 30204 711042
rect 29604 710722 29786 710958
rect 30022 710722 30204 710958
rect 26004 709438 26604 709460
rect 26004 709202 26186 709438
rect 26422 709202 26604 709438
rect 26004 709118 26604 709202
rect 26004 708882 26186 709118
rect 26422 708882 26604 709118
rect 22404 707598 23004 707620
rect 22404 707362 22586 707598
rect 22822 707362 23004 707598
rect 22404 707278 23004 707362
rect 22404 707042 22586 707278
rect 22822 707042 23004 707278
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7516 -6102 -7334 -5866
rect -7098 -6102 -6916 -5866
rect -7516 -6186 -6916 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 -6916 -6186
rect -7516 -6444 -6916 -6422
rect 11604 -5866 12204 12698
rect 18804 705758 19404 705780
rect 18804 705522 18986 705758
rect 19222 705522 19404 705758
rect 18804 705438 19404 705522
rect 18804 705202 18986 705438
rect 19222 705202 19404 705438
rect 18804 668454 19404 705202
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1266 19404 19898
rect 18804 -1502 18986 -1266
rect 19222 -1502 19404 -1266
rect 18804 -1586 19404 -1502
rect 18804 -1822 18986 -1586
rect 19222 -1822 19404 -1586
rect 18804 -1844 19404 -1822
rect 22404 672054 23004 707042
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3106 23004 23498
rect 22404 -3342 22586 -3106
rect 22822 -3342 23004 -3106
rect 22404 -3426 23004 -3342
rect 22404 -3662 22586 -3426
rect 22822 -3662 23004 -3426
rect 22404 -3684 23004 -3662
rect 26004 675654 26604 708882
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -4946 26604 27098
rect 26004 -5182 26186 -4946
rect 26422 -5182 26604 -4946
rect 26004 -5266 26604 -5182
rect 26004 -5502 26186 -5266
rect 26422 -5502 26604 -5266
rect 26004 -5524 26604 -5502
rect 29604 679254 30204 710722
rect 47604 710358 48204 711300
rect 47604 710122 47786 710358
rect 48022 710122 48204 710358
rect 47604 710038 48204 710122
rect 47604 709802 47786 710038
rect 48022 709802 48204 710038
rect 44004 708518 44604 709460
rect 44004 708282 44186 708518
rect 44422 708282 44604 708518
rect 44004 708198 44604 708282
rect 44004 707962 44186 708198
rect 44422 707962 44604 708198
rect 40404 706678 41004 707620
rect 40404 706442 40586 706678
rect 40822 706442 41004 706678
rect 40404 706358 41004 706442
rect 40404 706122 40586 706358
rect 40822 706122 41004 706358
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6102 11786 -5866
rect 12022 -6102 12204 -5866
rect 11604 -6186 12204 -6102
rect 11604 -6422 11786 -6186
rect 12022 -6422 12204 -6186
rect -8436 -7022 -8254 -6786
rect -8018 -7022 -7836 -6786
rect -8436 -7106 -7836 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 -7836 -7106
rect -8436 -7364 -7836 -7342
rect 11604 -7364 12204 -6422
rect 29604 -6786 30204 30698
rect 36804 704838 37404 705780
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1844 37404 -902
rect 40404 690054 41004 706122
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2186 41004 5498
rect 40404 -2422 40586 -2186
rect 40822 -2422 41004 -2186
rect 40404 -2506 41004 -2422
rect 40404 -2742 40586 -2506
rect 40822 -2742 41004 -2506
rect 40404 -3684 41004 -2742
rect 44004 693654 44604 707962
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4026 44604 9098
rect 44004 -4262 44186 -4026
rect 44422 -4262 44604 -4026
rect 44004 -4346 44604 -4262
rect 44004 -4582 44186 -4346
rect 44422 -4582 44604 -4346
rect 44004 -5524 44604 -4582
rect 47604 697254 48204 709802
rect 65604 711278 66204 711300
rect 65604 711042 65786 711278
rect 66022 711042 66204 711278
rect 65604 710958 66204 711042
rect 65604 710722 65786 710958
rect 66022 710722 66204 710958
rect 62004 709438 62604 709460
rect 62004 709202 62186 709438
rect 62422 709202 62604 709438
rect 62004 709118 62604 709202
rect 62004 708882 62186 709118
rect 62422 708882 62604 709118
rect 58404 707598 59004 707620
rect 58404 707362 58586 707598
rect 58822 707362 59004 707598
rect 58404 707278 59004 707362
rect 58404 707042 58586 707278
rect 58822 707042 59004 707278
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7022 29786 -6786
rect 30022 -7022 30204 -6786
rect 29604 -7106 30204 -7022
rect 29604 -7342 29786 -7106
rect 30022 -7342 30204 -7106
rect 29604 -7364 30204 -7342
rect 47604 -5866 48204 12698
rect 54804 705758 55404 705780
rect 54804 705522 54986 705758
rect 55222 705522 55404 705758
rect 54804 705438 55404 705522
rect 54804 705202 54986 705438
rect 55222 705202 55404 705438
rect 54804 668454 55404 705202
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1266 55404 19898
rect 54804 -1502 54986 -1266
rect 55222 -1502 55404 -1266
rect 54804 -1586 55404 -1502
rect 54804 -1822 54986 -1586
rect 55222 -1822 55404 -1586
rect 54804 -1844 55404 -1822
rect 58404 672054 59004 707042
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3106 59004 23498
rect 58404 -3342 58586 -3106
rect 58822 -3342 59004 -3106
rect 58404 -3426 59004 -3342
rect 58404 -3662 58586 -3426
rect 58822 -3662 59004 -3426
rect 58404 -3684 59004 -3662
rect 62004 675654 62604 708882
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 62004 531654 62604 567098
rect 62004 531418 62186 531654
rect 62422 531418 62604 531654
rect 62004 531334 62604 531418
rect 62004 531098 62186 531334
rect 62422 531098 62604 531334
rect 62004 495654 62604 531098
rect 62004 495418 62186 495654
rect 62422 495418 62604 495654
rect 62004 495334 62604 495418
rect 62004 495098 62186 495334
rect 62422 495098 62604 495334
rect 62004 459654 62604 495098
rect 62004 459418 62186 459654
rect 62422 459418 62604 459654
rect 62004 459334 62604 459418
rect 62004 459098 62186 459334
rect 62422 459098 62604 459334
rect 62004 423654 62604 459098
rect 62004 423418 62186 423654
rect 62422 423418 62604 423654
rect 62004 423334 62604 423418
rect 62004 423098 62186 423334
rect 62422 423098 62604 423334
rect 62004 387654 62604 423098
rect 62004 387418 62186 387654
rect 62422 387418 62604 387654
rect 62004 387334 62604 387418
rect 62004 387098 62186 387334
rect 62422 387098 62604 387334
rect 62004 351654 62604 387098
rect 62004 351418 62186 351654
rect 62422 351418 62604 351654
rect 62004 351334 62604 351418
rect 62004 351098 62186 351334
rect 62422 351098 62604 351334
rect 62004 315654 62604 351098
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -4946 62604 27098
rect 62004 -5182 62186 -4946
rect 62422 -5182 62604 -4946
rect 62004 -5266 62604 -5182
rect 62004 -5502 62186 -5266
rect 62422 -5502 62604 -5266
rect 62004 -5524 62604 -5502
rect 65604 679254 66204 710722
rect 83604 710358 84204 711300
rect 83604 710122 83786 710358
rect 84022 710122 84204 710358
rect 83604 710038 84204 710122
rect 83604 709802 83786 710038
rect 84022 709802 84204 710038
rect 80004 708518 80604 709460
rect 80004 708282 80186 708518
rect 80422 708282 80604 708518
rect 80004 708198 80604 708282
rect 80004 707962 80186 708198
rect 80422 707962 80604 708198
rect 76404 706678 77004 707620
rect 76404 706442 76586 706678
rect 76822 706442 77004 706678
rect 76404 706358 77004 706442
rect 76404 706122 76586 706358
rect 76822 706122 77004 706358
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 65604 571254 66204 606698
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 535254 66204 570698
rect 65604 535018 65786 535254
rect 66022 535018 66204 535254
rect 65604 534934 66204 535018
rect 65604 534698 65786 534934
rect 66022 534698 66204 534934
rect 65604 499254 66204 534698
rect 65604 499018 65786 499254
rect 66022 499018 66204 499254
rect 65604 498934 66204 499018
rect 65604 498698 65786 498934
rect 66022 498698 66204 498934
rect 65604 463254 66204 498698
rect 65604 463018 65786 463254
rect 66022 463018 66204 463254
rect 65604 462934 66204 463018
rect 65604 462698 65786 462934
rect 66022 462698 66204 462934
rect 65604 427254 66204 462698
rect 65604 427018 65786 427254
rect 66022 427018 66204 427254
rect 65604 426934 66204 427018
rect 65604 426698 65786 426934
rect 66022 426698 66204 426934
rect 65604 391254 66204 426698
rect 65604 391018 65786 391254
rect 66022 391018 66204 391254
rect 65604 390934 66204 391018
rect 65604 390698 65786 390934
rect 66022 390698 66204 390934
rect 65604 355254 66204 390698
rect 65604 355018 65786 355254
rect 66022 355018 66204 355254
rect 65604 354934 66204 355018
rect 65604 354698 65786 354934
rect 66022 354698 66204 354934
rect 65604 319254 66204 354698
rect 65604 319018 65786 319254
rect 66022 319018 66204 319254
rect 65604 318934 66204 319018
rect 65604 318698 65786 318934
rect 66022 318698 66204 318934
rect 65604 283254 66204 318698
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6102 47786 -5866
rect 48022 -6102 48204 -5866
rect 47604 -6186 48204 -6102
rect 47604 -6422 47786 -6186
rect 48022 -6422 48204 -6186
rect 47604 -7364 48204 -6422
rect 65604 -6786 66204 30698
rect 72804 704838 73404 705780
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1844 73404 -902
rect 76404 690054 77004 706122
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 366054 77004 401498
rect 76404 365818 76586 366054
rect 76822 365818 77004 366054
rect 76404 365734 77004 365818
rect 76404 365498 76586 365734
rect 76822 365498 77004 365734
rect 76404 330054 77004 365498
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2186 77004 5498
rect 76404 -2422 76586 -2186
rect 76822 -2422 77004 -2186
rect 76404 -2506 77004 -2422
rect 76404 -2742 76586 -2506
rect 76822 -2742 77004 -2506
rect 76404 -3684 77004 -2742
rect 80004 693654 80604 707962
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 621654 80604 657098
rect 80004 621418 80186 621654
rect 80422 621418 80604 621654
rect 80004 621334 80604 621418
rect 80004 621098 80186 621334
rect 80422 621098 80604 621334
rect 80004 585654 80604 621098
rect 80004 585418 80186 585654
rect 80422 585418 80604 585654
rect 80004 585334 80604 585418
rect 80004 585098 80186 585334
rect 80422 585098 80604 585334
rect 80004 549654 80604 585098
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 513654 80604 549098
rect 80004 513418 80186 513654
rect 80422 513418 80604 513654
rect 80004 513334 80604 513418
rect 80004 513098 80186 513334
rect 80422 513098 80604 513334
rect 80004 477654 80604 513098
rect 80004 477418 80186 477654
rect 80422 477418 80604 477654
rect 80004 477334 80604 477418
rect 80004 477098 80186 477334
rect 80422 477098 80604 477334
rect 80004 441654 80604 477098
rect 80004 441418 80186 441654
rect 80422 441418 80604 441654
rect 80004 441334 80604 441418
rect 80004 441098 80186 441334
rect 80422 441098 80604 441334
rect 80004 405654 80604 441098
rect 80004 405418 80186 405654
rect 80422 405418 80604 405654
rect 80004 405334 80604 405418
rect 80004 405098 80186 405334
rect 80422 405098 80604 405334
rect 80004 369654 80604 405098
rect 80004 369418 80186 369654
rect 80422 369418 80604 369654
rect 80004 369334 80604 369418
rect 80004 369098 80186 369334
rect 80422 369098 80604 369334
rect 80004 333654 80604 369098
rect 80004 333418 80186 333654
rect 80422 333418 80604 333654
rect 80004 333334 80604 333418
rect 80004 333098 80186 333334
rect 80422 333098 80604 333334
rect 80004 297654 80604 333098
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4026 80604 9098
rect 80004 -4262 80186 -4026
rect 80422 -4262 80604 -4026
rect 80004 -4346 80604 -4262
rect 80004 -4582 80186 -4346
rect 80422 -4582 80604 -4346
rect 80004 -5524 80604 -4582
rect 83604 697254 84204 709802
rect 101604 711278 102204 711300
rect 101604 711042 101786 711278
rect 102022 711042 102204 711278
rect 101604 710958 102204 711042
rect 101604 710722 101786 710958
rect 102022 710722 102204 710958
rect 98004 709438 98604 709460
rect 98004 709202 98186 709438
rect 98422 709202 98604 709438
rect 98004 709118 98604 709202
rect 98004 708882 98186 709118
rect 98422 708882 98604 709118
rect 94404 707598 95004 707620
rect 94404 707362 94586 707598
rect 94822 707362 95004 707598
rect 94404 707278 95004 707362
rect 94404 707042 94586 707278
rect 94822 707042 95004 707278
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 625254 84204 660698
rect 83604 625018 83786 625254
rect 84022 625018 84204 625254
rect 83604 624934 84204 625018
rect 83604 624698 83786 624934
rect 84022 624698 84204 624934
rect 83604 589254 84204 624698
rect 83604 589018 83786 589254
rect 84022 589018 84204 589254
rect 83604 588934 84204 589018
rect 83604 588698 83786 588934
rect 84022 588698 84204 588934
rect 83604 553254 84204 588698
rect 83604 553018 83786 553254
rect 84022 553018 84204 553254
rect 83604 552934 84204 553018
rect 83604 552698 83786 552934
rect 84022 552698 84204 552934
rect 83604 517254 84204 552698
rect 83604 517018 83786 517254
rect 84022 517018 84204 517254
rect 83604 516934 84204 517018
rect 83604 516698 83786 516934
rect 84022 516698 84204 516934
rect 83604 481254 84204 516698
rect 83604 481018 83786 481254
rect 84022 481018 84204 481254
rect 83604 480934 84204 481018
rect 83604 480698 83786 480934
rect 84022 480698 84204 480934
rect 83604 445254 84204 480698
rect 83604 445018 83786 445254
rect 84022 445018 84204 445254
rect 83604 444934 84204 445018
rect 83604 444698 83786 444934
rect 84022 444698 84204 444934
rect 83604 409254 84204 444698
rect 83604 409018 83786 409254
rect 84022 409018 84204 409254
rect 83604 408934 84204 409018
rect 83604 408698 83786 408934
rect 84022 408698 84204 408934
rect 83604 373254 84204 408698
rect 83604 373018 83786 373254
rect 84022 373018 84204 373254
rect 83604 372934 84204 373018
rect 83604 372698 83786 372934
rect 84022 372698 84204 372934
rect 83604 337254 84204 372698
rect 83604 337018 83786 337254
rect 84022 337018 84204 337254
rect 83604 336934 84204 337018
rect 83604 336698 83786 336934
rect 84022 336698 84204 336934
rect 83604 301254 84204 336698
rect 83604 301018 83786 301254
rect 84022 301018 84204 301254
rect 83604 300934 84204 301018
rect 83604 300698 83786 300934
rect 84022 300698 84204 300934
rect 83604 265254 84204 300698
rect 83604 265018 83786 265254
rect 84022 265018 84204 265254
rect 83604 264934 84204 265018
rect 83604 264698 83786 264934
rect 84022 264698 84204 264934
rect 83604 229254 84204 264698
rect 83604 229018 83786 229254
rect 84022 229018 84204 229254
rect 83604 228934 84204 229018
rect 83604 228698 83786 228934
rect 84022 228698 84204 228934
rect 83604 193254 84204 228698
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7022 65786 -6786
rect 66022 -7022 66204 -6786
rect 65604 -7106 66204 -7022
rect 65604 -7342 65786 -7106
rect 66022 -7342 66204 -7106
rect 65604 -7364 66204 -7342
rect 83604 -5866 84204 12698
rect 90804 705758 91404 705780
rect 90804 705522 90986 705758
rect 91222 705522 91404 705758
rect 90804 705438 91404 705522
rect 90804 705202 90986 705438
rect 91222 705202 91404 705438
rect 90804 668454 91404 705202
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 560454 91404 595898
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 524454 91404 559898
rect 90804 524218 90986 524454
rect 91222 524218 91404 524454
rect 90804 524134 91404 524218
rect 90804 523898 90986 524134
rect 91222 523898 91404 524134
rect 90804 488454 91404 523898
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 452454 91404 487898
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 416454 91404 451898
rect 90804 416218 90986 416454
rect 91222 416218 91404 416454
rect 90804 416134 91404 416218
rect 90804 415898 90986 416134
rect 91222 415898 91404 416134
rect 90804 380454 91404 415898
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 90804 344454 91404 379898
rect 90804 344218 90986 344454
rect 91222 344218 91404 344454
rect 90804 344134 91404 344218
rect 90804 343898 90986 344134
rect 91222 343898 91404 344134
rect 90804 308454 91404 343898
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1266 91404 19898
rect 90804 -1502 90986 -1266
rect 91222 -1502 91404 -1266
rect 90804 -1586 91404 -1502
rect 90804 -1822 90986 -1586
rect 91222 -1822 91404 -1586
rect 90804 -1844 91404 -1822
rect 94404 672054 95004 707042
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 600054 95004 635498
rect 94404 599818 94586 600054
rect 94822 599818 95004 600054
rect 94404 599734 95004 599818
rect 94404 599498 94586 599734
rect 94822 599498 95004 599734
rect 94404 564054 95004 599498
rect 94404 563818 94586 564054
rect 94822 563818 95004 564054
rect 94404 563734 95004 563818
rect 94404 563498 94586 563734
rect 94822 563498 95004 563734
rect 94404 528054 95004 563498
rect 94404 527818 94586 528054
rect 94822 527818 95004 528054
rect 94404 527734 95004 527818
rect 94404 527498 94586 527734
rect 94822 527498 95004 527734
rect 94404 492054 95004 527498
rect 94404 491818 94586 492054
rect 94822 491818 95004 492054
rect 94404 491734 95004 491818
rect 94404 491498 94586 491734
rect 94822 491498 95004 491734
rect 94404 456054 95004 491498
rect 94404 455818 94586 456054
rect 94822 455818 95004 456054
rect 94404 455734 95004 455818
rect 94404 455498 94586 455734
rect 94822 455498 95004 455734
rect 94404 420054 95004 455498
rect 94404 419818 94586 420054
rect 94822 419818 95004 420054
rect 94404 419734 95004 419818
rect 94404 419498 94586 419734
rect 94822 419498 95004 419734
rect 94404 384054 95004 419498
rect 94404 383818 94586 384054
rect 94822 383818 95004 384054
rect 94404 383734 95004 383818
rect 94404 383498 94586 383734
rect 94822 383498 95004 383734
rect 94404 348054 95004 383498
rect 94404 347818 94586 348054
rect 94822 347818 95004 348054
rect 94404 347734 95004 347818
rect 94404 347498 94586 347734
rect 94822 347498 95004 347734
rect 94404 312054 95004 347498
rect 94404 311818 94586 312054
rect 94822 311818 95004 312054
rect 94404 311734 95004 311818
rect 94404 311498 94586 311734
rect 94822 311498 95004 311734
rect 94404 276054 95004 311498
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3106 95004 23498
rect 94404 -3342 94586 -3106
rect 94822 -3342 95004 -3106
rect 94404 -3426 95004 -3342
rect 94404 -3662 94586 -3426
rect 94822 -3662 95004 -3426
rect 94404 -3684 95004 -3662
rect 98004 675654 98604 708882
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 639654 98604 675098
rect 98004 639418 98186 639654
rect 98422 639418 98604 639654
rect 98004 639334 98604 639418
rect 98004 639098 98186 639334
rect 98422 639098 98604 639334
rect 98004 603654 98604 639098
rect 98004 603418 98186 603654
rect 98422 603418 98604 603654
rect 98004 603334 98604 603418
rect 98004 603098 98186 603334
rect 98422 603098 98604 603334
rect 98004 567654 98604 603098
rect 98004 567418 98186 567654
rect 98422 567418 98604 567654
rect 98004 567334 98604 567418
rect 98004 567098 98186 567334
rect 98422 567098 98604 567334
rect 98004 531654 98604 567098
rect 98004 531418 98186 531654
rect 98422 531418 98604 531654
rect 98004 531334 98604 531418
rect 98004 531098 98186 531334
rect 98422 531098 98604 531334
rect 98004 495654 98604 531098
rect 98004 495418 98186 495654
rect 98422 495418 98604 495654
rect 98004 495334 98604 495418
rect 98004 495098 98186 495334
rect 98422 495098 98604 495334
rect 98004 459654 98604 495098
rect 98004 459418 98186 459654
rect 98422 459418 98604 459654
rect 98004 459334 98604 459418
rect 98004 459098 98186 459334
rect 98422 459098 98604 459334
rect 98004 423654 98604 459098
rect 98004 423418 98186 423654
rect 98422 423418 98604 423654
rect 98004 423334 98604 423418
rect 98004 423098 98186 423334
rect 98422 423098 98604 423334
rect 98004 387654 98604 423098
rect 98004 387418 98186 387654
rect 98422 387418 98604 387654
rect 98004 387334 98604 387418
rect 98004 387098 98186 387334
rect 98422 387098 98604 387334
rect 98004 351654 98604 387098
rect 98004 351418 98186 351654
rect 98422 351418 98604 351654
rect 98004 351334 98604 351418
rect 98004 351098 98186 351334
rect 98422 351098 98604 351334
rect 98004 315654 98604 351098
rect 98004 315418 98186 315654
rect 98422 315418 98604 315654
rect 98004 315334 98604 315418
rect 98004 315098 98186 315334
rect 98422 315098 98604 315334
rect 98004 279654 98604 315098
rect 98004 279418 98186 279654
rect 98422 279418 98604 279654
rect 98004 279334 98604 279418
rect 98004 279098 98186 279334
rect 98422 279098 98604 279334
rect 98004 243654 98604 279098
rect 98004 243418 98186 243654
rect 98422 243418 98604 243654
rect 98004 243334 98604 243418
rect 98004 243098 98186 243334
rect 98422 243098 98604 243334
rect 98004 207654 98604 243098
rect 98004 207418 98186 207654
rect 98422 207418 98604 207654
rect 98004 207334 98604 207418
rect 98004 207098 98186 207334
rect 98422 207098 98604 207334
rect 98004 171654 98604 207098
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -4946 98604 27098
rect 98004 -5182 98186 -4946
rect 98422 -5182 98604 -4946
rect 98004 -5266 98604 -5182
rect 98004 -5502 98186 -5266
rect 98422 -5502 98604 -5266
rect 98004 -5524 98604 -5502
rect 101604 679254 102204 710722
rect 119604 710358 120204 711300
rect 119604 710122 119786 710358
rect 120022 710122 120204 710358
rect 119604 710038 120204 710122
rect 119604 709802 119786 710038
rect 120022 709802 120204 710038
rect 116004 708518 116604 709460
rect 116004 708282 116186 708518
rect 116422 708282 116604 708518
rect 116004 708198 116604 708282
rect 116004 707962 116186 708198
rect 116422 707962 116604 708198
rect 112404 706678 113004 707620
rect 112404 706442 112586 706678
rect 112822 706442 113004 706678
rect 112404 706358 113004 706442
rect 112404 706122 112586 706358
rect 112822 706122 113004 706358
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 643254 102204 678698
rect 101604 643018 101786 643254
rect 102022 643018 102204 643254
rect 101604 642934 102204 643018
rect 101604 642698 101786 642934
rect 102022 642698 102204 642934
rect 101604 607254 102204 642698
rect 101604 607018 101786 607254
rect 102022 607018 102204 607254
rect 101604 606934 102204 607018
rect 101604 606698 101786 606934
rect 102022 606698 102204 606934
rect 101604 571254 102204 606698
rect 101604 571018 101786 571254
rect 102022 571018 102204 571254
rect 101604 570934 102204 571018
rect 101604 570698 101786 570934
rect 102022 570698 102204 570934
rect 101604 535254 102204 570698
rect 101604 535018 101786 535254
rect 102022 535018 102204 535254
rect 101604 534934 102204 535018
rect 101604 534698 101786 534934
rect 102022 534698 102204 534934
rect 101604 499254 102204 534698
rect 101604 499018 101786 499254
rect 102022 499018 102204 499254
rect 101604 498934 102204 499018
rect 101604 498698 101786 498934
rect 102022 498698 102204 498934
rect 101604 463254 102204 498698
rect 101604 463018 101786 463254
rect 102022 463018 102204 463254
rect 101604 462934 102204 463018
rect 101604 462698 101786 462934
rect 102022 462698 102204 462934
rect 101604 427254 102204 462698
rect 101604 427018 101786 427254
rect 102022 427018 102204 427254
rect 101604 426934 102204 427018
rect 101604 426698 101786 426934
rect 102022 426698 102204 426934
rect 101604 391254 102204 426698
rect 101604 391018 101786 391254
rect 102022 391018 102204 391254
rect 101604 390934 102204 391018
rect 101604 390698 101786 390934
rect 102022 390698 102204 390934
rect 101604 355254 102204 390698
rect 101604 355018 101786 355254
rect 102022 355018 102204 355254
rect 101604 354934 102204 355018
rect 101604 354698 101786 354934
rect 102022 354698 102204 354934
rect 101604 319254 102204 354698
rect 101604 319018 101786 319254
rect 102022 319018 102204 319254
rect 101604 318934 102204 319018
rect 101604 318698 101786 318934
rect 102022 318698 102204 318934
rect 101604 283254 102204 318698
rect 101604 283018 101786 283254
rect 102022 283018 102204 283254
rect 101604 282934 102204 283018
rect 101604 282698 101786 282934
rect 102022 282698 102204 282934
rect 101604 247254 102204 282698
rect 101604 247018 101786 247254
rect 102022 247018 102204 247254
rect 101604 246934 102204 247018
rect 101604 246698 101786 246934
rect 102022 246698 102204 246934
rect 101604 211254 102204 246698
rect 101604 211018 101786 211254
rect 102022 211018 102204 211254
rect 101604 210934 102204 211018
rect 101604 210698 101786 210934
rect 102022 210698 102204 210934
rect 101604 175254 102204 210698
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6102 83786 -5866
rect 84022 -6102 84204 -5866
rect 83604 -6186 84204 -6102
rect 83604 -6422 83786 -6186
rect 84022 -6422 84204 -6186
rect 83604 -7364 84204 -6422
rect 101604 -6786 102204 30698
rect 108804 704838 109404 705780
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 578454 109404 613898
rect 108804 578218 108986 578454
rect 109222 578218 109404 578454
rect 108804 578134 109404 578218
rect 108804 577898 108986 578134
rect 109222 577898 109404 578134
rect 108804 542454 109404 577898
rect 108804 542218 108986 542454
rect 109222 542218 109404 542454
rect 108804 542134 109404 542218
rect 108804 541898 108986 542134
rect 109222 541898 109404 542134
rect 108804 506454 109404 541898
rect 108804 506218 108986 506454
rect 109222 506218 109404 506454
rect 108804 506134 109404 506218
rect 108804 505898 108986 506134
rect 109222 505898 109404 506134
rect 108804 470454 109404 505898
rect 108804 470218 108986 470454
rect 109222 470218 109404 470454
rect 108804 470134 109404 470218
rect 108804 469898 108986 470134
rect 109222 469898 109404 470134
rect 108804 434454 109404 469898
rect 108804 434218 108986 434454
rect 109222 434218 109404 434454
rect 108804 434134 109404 434218
rect 108804 433898 108986 434134
rect 109222 433898 109404 434134
rect 108804 398454 109404 433898
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 362454 109404 397898
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 326454 109404 361898
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1844 109404 -902
rect 112404 690054 113004 706122
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 582054 113004 617498
rect 112404 581818 112586 582054
rect 112822 581818 113004 582054
rect 112404 581734 113004 581818
rect 112404 581498 112586 581734
rect 112822 581498 113004 581734
rect 112404 546054 113004 581498
rect 112404 545818 112586 546054
rect 112822 545818 113004 546054
rect 112404 545734 113004 545818
rect 112404 545498 112586 545734
rect 112822 545498 113004 545734
rect 112404 510054 113004 545498
rect 112404 509818 112586 510054
rect 112822 509818 113004 510054
rect 112404 509734 113004 509818
rect 112404 509498 112586 509734
rect 112822 509498 113004 509734
rect 112404 474054 113004 509498
rect 112404 473818 112586 474054
rect 112822 473818 113004 474054
rect 112404 473734 113004 473818
rect 112404 473498 112586 473734
rect 112822 473498 113004 473734
rect 112404 438054 113004 473498
rect 112404 437818 112586 438054
rect 112822 437818 113004 438054
rect 112404 437734 113004 437818
rect 112404 437498 112586 437734
rect 112822 437498 113004 437734
rect 112404 402054 113004 437498
rect 112404 401818 112586 402054
rect 112822 401818 113004 402054
rect 112404 401734 113004 401818
rect 112404 401498 112586 401734
rect 112822 401498 113004 401734
rect 112404 366054 113004 401498
rect 112404 365818 112586 366054
rect 112822 365818 113004 366054
rect 112404 365734 113004 365818
rect 112404 365498 112586 365734
rect 112822 365498 113004 365734
rect 112404 330054 113004 365498
rect 112404 329818 112586 330054
rect 112822 329818 113004 330054
rect 112404 329734 113004 329818
rect 112404 329498 112586 329734
rect 112822 329498 113004 329734
rect 112404 294054 113004 329498
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2186 113004 5498
rect 112404 -2422 112586 -2186
rect 112822 -2422 113004 -2186
rect 112404 -2506 113004 -2422
rect 112404 -2742 112586 -2506
rect 112822 -2742 113004 -2506
rect 112404 -3684 113004 -2742
rect 116004 693654 116604 707962
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 621654 116604 657098
rect 116004 621418 116186 621654
rect 116422 621418 116604 621654
rect 116004 621334 116604 621418
rect 116004 621098 116186 621334
rect 116422 621098 116604 621334
rect 116004 585654 116604 621098
rect 116004 585418 116186 585654
rect 116422 585418 116604 585654
rect 116004 585334 116604 585418
rect 116004 585098 116186 585334
rect 116422 585098 116604 585334
rect 116004 549654 116604 585098
rect 116004 549418 116186 549654
rect 116422 549418 116604 549654
rect 116004 549334 116604 549418
rect 116004 549098 116186 549334
rect 116422 549098 116604 549334
rect 116004 513654 116604 549098
rect 116004 513418 116186 513654
rect 116422 513418 116604 513654
rect 116004 513334 116604 513418
rect 116004 513098 116186 513334
rect 116422 513098 116604 513334
rect 116004 477654 116604 513098
rect 116004 477418 116186 477654
rect 116422 477418 116604 477654
rect 116004 477334 116604 477418
rect 116004 477098 116186 477334
rect 116422 477098 116604 477334
rect 116004 441654 116604 477098
rect 116004 441418 116186 441654
rect 116422 441418 116604 441654
rect 116004 441334 116604 441418
rect 116004 441098 116186 441334
rect 116422 441098 116604 441334
rect 116004 405654 116604 441098
rect 116004 405418 116186 405654
rect 116422 405418 116604 405654
rect 116004 405334 116604 405418
rect 116004 405098 116186 405334
rect 116422 405098 116604 405334
rect 116004 369654 116604 405098
rect 116004 369418 116186 369654
rect 116422 369418 116604 369654
rect 116004 369334 116604 369418
rect 116004 369098 116186 369334
rect 116422 369098 116604 369334
rect 116004 333654 116604 369098
rect 116004 333418 116186 333654
rect 116422 333418 116604 333654
rect 116004 333334 116604 333418
rect 116004 333098 116186 333334
rect 116422 333098 116604 333334
rect 116004 297654 116604 333098
rect 116004 297418 116186 297654
rect 116422 297418 116604 297654
rect 116004 297334 116604 297418
rect 116004 297098 116186 297334
rect 116422 297098 116604 297334
rect 116004 261654 116604 297098
rect 116004 261418 116186 261654
rect 116422 261418 116604 261654
rect 116004 261334 116604 261418
rect 116004 261098 116186 261334
rect 116422 261098 116604 261334
rect 116004 225654 116604 261098
rect 116004 225418 116186 225654
rect 116422 225418 116604 225654
rect 116004 225334 116604 225418
rect 116004 225098 116186 225334
rect 116422 225098 116604 225334
rect 116004 189654 116604 225098
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4026 116604 9098
rect 116004 -4262 116186 -4026
rect 116422 -4262 116604 -4026
rect 116004 -4346 116604 -4262
rect 116004 -4582 116186 -4346
rect 116422 -4582 116604 -4346
rect 116004 -5524 116604 -4582
rect 119604 697254 120204 709802
rect 137604 711278 138204 711300
rect 137604 711042 137786 711278
rect 138022 711042 138204 711278
rect 137604 710958 138204 711042
rect 137604 710722 137786 710958
rect 138022 710722 138204 710958
rect 134004 709438 134604 709460
rect 134004 709202 134186 709438
rect 134422 709202 134604 709438
rect 134004 709118 134604 709202
rect 134004 708882 134186 709118
rect 134422 708882 134604 709118
rect 130404 707598 131004 707620
rect 130404 707362 130586 707598
rect 130822 707362 131004 707598
rect 130404 707278 131004 707362
rect 130404 707042 130586 707278
rect 130822 707042 131004 707278
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 625254 120204 660698
rect 119604 625018 119786 625254
rect 120022 625018 120204 625254
rect 119604 624934 120204 625018
rect 119604 624698 119786 624934
rect 120022 624698 120204 624934
rect 119604 589254 120204 624698
rect 119604 589018 119786 589254
rect 120022 589018 120204 589254
rect 119604 588934 120204 589018
rect 119604 588698 119786 588934
rect 120022 588698 120204 588934
rect 119604 553254 120204 588698
rect 119604 553018 119786 553254
rect 120022 553018 120204 553254
rect 119604 552934 120204 553018
rect 119604 552698 119786 552934
rect 120022 552698 120204 552934
rect 119604 517254 120204 552698
rect 119604 517018 119786 517254
rect 120022 517018 120204 517254
rect 119604 516934 120204 517018
rect 119604 516698 119786 516934
rect 120022 516698 120204 516934
rect 119604 481254 120204 516698
rect 119604 481018 119786 481254
rect 120022 481018 120204 481254
rect 119604 480934 120204 481018
rect 119604 480698 119786 480934
rect 120022 480698 120204 480934
rect 119604 445254 120204 480698
rect 119604 445018 119786 445254
rect 120022 445018 120204 445254
rect 119604 444934 120204 445018
rect 119604 444698 119786 444934
rect 120022 444698 120204 444934
rect 119604 409254 120204 444698
rect 119604 409018 119786 409254
rect 120022 409018 120204 409254
rect 119604 408934 120204 409018
rect 119604 408698 119786 408934
rect 120022 408698 120204 408934
rect 119604 373254 120204 408698
rect 119604 373018 119786 373254
rect 120022 373018 120204 373254
rect 119604 372934 120204 373018
rect 119604 372698 119786 372934
rect 120022 372698 120204 372934
rect 119604 337254 120204 372698
rect 119604 337018 119786 337254
rect 120022 337018 120204 337254
rect 119604 336934 120204 337018
rect 119604 336698 119786 336934
rect 120022 336698 120204 336934
rect 119604 301254 120204 336698
rect 119604 301018 119786 301254
rect 120022 301018 120204 301254
rect 119604 300934 120204 301018
rect 119604 300698 119786 300934
rect 120022 300698 120204 300934
rect 119604 265254 120204 300698
rect 119604 265018 119786 265254
rect 120022 265018 120204 265254
rect 119604 264934 120204 265018
rect 119604 264698 119786 264934
rect 120022 264698 120204 264934
rect 119604 229254 120204 264698
rect 119604 229018 119786 229254
rect 120022 229018 120204 229254
rect 119604 228934 120204 229018
rect 119604 228698 119786 228934
rect 120022 228698 120204 228934
rect 119604 193254 120204 228698
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7022 101786 -6786
rect 102022 -7022 102204 -6786
rect 101604 -7106 102204 -7022
rect 101604 -7342 101786 -7106
rect 102022 -7342 102204 -7106
rect 101604 -7364 102204 -7342
rect 119604 -5866 120204 12698
rect 126804 705758 127404 705780
rect 126804 705522 126986 705758
rect 127222 705522 127404 705758
rect 126804 705438 127404 705522
rect 126804 705202 126986 705438
rect 127222 705202 127404 705438
rect 126804 668454 127404 705202
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 560454 127404 595898
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 524454 127404 559898
rect 126804 524218 126986 524454
rect 127222 524218 127404 524454
rect 126804 524134 127404 524218
rect 126804 523898 126986 524134
rect 127222 523898 127404 524134
rect 126804 488454 127404 523898
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 452454 127404 487898
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 416454 127404 451898
rect 126804 416218 126986 416454
rect 127222 416218 127404 416454
rect 126804 416134 127404 416218
rect 126804 415898 126986 416134
rect 127222 415898 127404 416134
rect 126804 380454 127404 415898
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1266 127404 19898
rect 126804 -1502 126986 -1266
rect 127222 -1502 127404 -1266
rect 126804 -1586 127404 -1502
rect 126804 -1822 126986 -1586
rect 127222 -1822 127404 -1586
rect 126804 -1844 127404 -1822
rect 130404 672054 131004 707042
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 600054 131004 635498
rect 130404 599818 130586 600054
rect 130822 599818 131004 600054
rect 130404 599734 131004 599818
rect 130404 599498 130586 599734
rect 130822 599498 131004 599734
rect 130404 564054 131004 599498
rect 130404 563818 130586 564054
rect 130822 563818 131004 564054
rect 130404 563734 131004 563818
rect 130404 563498 130586 563734
rect 130822 563498 131004 563734
rect 130404 528054 131004 563498
rect 130404 527818 130586 528054
rect 130822 527818 131004 528054
rect 130404 527734 131004 527818
rect 130404 527498 130586 527734
rect 130822 527498 131004 527734
rect 130404 492054 131004 527498
rect 130404 491818 130586 492054
rect 130822 491818 131004 492054
rect 130404 491734 131004 491818
rect 130404 491498 130586 491734
rect 130822 491498 131004 491734
rect 130404 456054 131004 491498
rect 130404 455818 130586 456054
rect 130822 455818 131004 456054
rect 130404 455734 131004 455818
rect 130404 455498 130586 455734
rect 130822 455498 131004 455734
rect 130404 420054 131004 455498
rect 130404 419818 130586 420054
rect 130822 419818 131004 420054
rect 130404 419734 131004 419818
rect 130404 419498 130586 419734
rect 130822 419498 131004 419734
rect 130404 384054 131004 419498
rect 130404 383818 130586 384054
rect 130822 383818 131004 384054
rect 130404 383734 131004 383818
rect 130404 383498 130586 383734
rect 130822 383498 131004 383734
rect 130404 348054 131004 383498
rect 130404 347818 130586 348054
rect 130822 347818 131004 348054
rect 130404 347734 131004 347818
rect 130404 347498 130586 347734
rect 130822 347498 131004 347734
rect 130404 312054 131004 347498
rect 130404 311818 130586 312054
rect 130822 311818 131004 312054
rect 130404 311734 131004 311818
rect 130404 311498 130586 311734
rect 130822 311498 131004 311734
rect 130404 276054 131004 311498
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3106 131004 23498
rect 130404 -3342 130586 -3106
rect 130822 -3342 131004 -3106
rect 130404 -3426 131004 -3342
rect 130404 -3662 130586 -3426
rect 130822 -3662 131004 -3426
rect 130404 -3684 131004 -3662
rect 134004 675654 134604 708882
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 639654 134604 675098
rect 134004 639418 134186 639654
rect 134422 639418 134604 639654
rect 134004 639334 134604 639418
rect 134004 639098 134186 639334
rect 134422 639098 134604 639334
rect 134004 603654 134604 639098
rect 134004 603418 134186 603654
rect 134422 603418 134604 603654
rect 134004 603334 134604 603418
rect 134004 603098 134186 603334
rect 134422 603098 134604 603334
rect 134004 567654 134604 603098
rect 134004 567418 134186 567654
rect 134422 567418 134604 567654
rect 134004 567334 134604 567418
rect 134004 567098 134186 567334
rect 134422 567098 134604 567334
rect 134004 531654 134604 567098
rect 134004 531418 134186 531654
rect 134422 531418 134604 531654
rect 134004 531334 134604 531418
rect 134004 531098 134186 531334
rect 134422 531098 134604 531334
rect 134004 495654 134604 531098
rect 134004 495418 134186 495654
rect 134422 495418 134604 495654
rect 134004 495334 134604 495418
rect 134004 495098 134186 495334
rect 134422 495098 134604 495334
rect 134004 459654 134604 495098
rect 134004 459418 134186 459654
rect 134422 459418 134604 459654
rect 134004 459334 134604 459418
rect 134004 459098 134186 459334
rect 134422 459098 134604 459334
rect 134004 423654 134604 459098
rect 134004 423418 134186 423654
rect 134422 423418 134604 423654
rect 134004 423334 134604 423418
rect 134004 423098 134186 423334
rect 134422 423098 134604 423334
rect 134004 387654 134604 423098
rect 134004 387418 134186 387654
rect 134422 387418 134604 387654
rect 134004 387334 134604 387418
rect 134004 387098 134186 387334
rect 134422 387098 134604 387334
rect 134004 351654 134604 387098
rect 134004 351418 134186 351654
rect 134422 351418 134604 351654
rect 134004 351334 134604 351418
rect 134004 351098 134186 351334
rect 134422 351098 134604 351334
rect 134004 315654 134604 351098
rect 134004 315418 134186 315654
rect 134422 315418 134604 315654
rect 134004 315334 134604 315418
rect 134004 315098 134186 315334
rect 134422 315098 134604 315334
rect 134004 279654 134604 315098
rect 134004 279418 134186 279654
rect 134422 279418 134604 279654
rect 134004 279334 134604 279418
rect 134004 279098 134186 279334
rect 134422 279098 134604 279334
rect 134004 243654 134604 279098
rect 134004 243418 134186 243654
rect 134422 243418 134604 243654
rect 134004 243334 134604 243418
rect 134004 243098 134186 243334
rect 134422 243098 134604 243334
rect 134004 207654 134604 243098
rect 134004 207418 134186 207654
rect 134422 207418 134604 207654
rect 134004 207334 134604 207418
rect 134004 207098 134186 207334
rect 134422 207098 134604 207334
rect 134004 171654 134604 207098
rect 134004 171418 134186 171654
rect 134422 171418 134604 171654
rect 134004 171334 134604 171418
rect 134004 171098 134186 171334
rect 134422 171098 134604 171334
rect 134004 135654 134604 171098
rect 134004 135418 134186 135654
rect 134422 135418 134604 135654
rect 134004 135334 134604 135418
rect 134004 135098 134186 135334
rect 134422 135098 134604 135334
rect 134004 99654 134604 135098
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -4946 134604 27098
rect 134004 -5182 134186 -4946
rect 134422 -5182 134604 -4946
rect 134004 -5266 134604 -5182
rect 134004 -5502 134186 -5266
rect 134422 -5502 134604 -5266
rect 134004 -5524 134604 -5502
rect 137604 679254 138204 710722
rect 155604 710358 156204 711300
rect 155604 710122 155786 710358
rect 156022 710122 156204 710358
rect 155604 710038 156204 710122
rect 155604 709802 155786 710038
rect 156022 709802 156204 710038
rect 152004 708518 152604 709460
rect 152004 708282 152186 708518
rect 152422 708282 152604 708518
rect 152004 708198 152604 708282
rect 152004 707962 152186 708198
rect 152422 707962 152604 708198
rect 148404 706678 149004 707620
rect 148404 706442 148586 706678
rect 148822 706442 149004 706678
rect 148404 706358 149004 706442
rect 148404 706122 148586 706358
rect 148822 706122 149004 706358
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 643254 138204 678698
rect 137604 643018 137786 643254
rect 138022 643018 138204 643254
rect 137604 642934 138204 643018
rect 137604 642698 137786 642934
rect 138022 642698 138204 642934
rect 137604 607254 138204 642698
rect 137604 607018 137786 607254
rect 138022 607018 138204 607254
rect 137604 606934 138204 607018
rect 137604 606698 137786 606934
rect 138022 606698 138204 606934
rect 137604 571254 138204 606698
rect 137604 571018 137786 571254
rect 138022 571018 138204 571254
rect 137604 570934 138204 571018
rect 137604 570698 137786 570934
rect 138022 570698 138204 570934
rect 137604 535254 138204 570698
rect 137604 535018 137786 535254
rect 138022 535018 138204 535254
rect 137604 534934 138204 535018
rect 137604 534698 137786 534934
rect 138022 534698 138204 534934
rect 137604 499254 138204 534698
rect 137604 499018 137786 499254
rect 138022 499018 138204 499254
rect 137604 498934 138204 499018
rect 137604 498698 137786 498934
rect 138022 498698 138204 498934
rect 137604 463254 138204 498698
rect 137604 463018 137786 463254
rect 138022 463018 138204 463254
rect 137604 462934 138204 463018
rect 137604 462698 137786 462934
rect 138022 462698 138204 462934
rect 137604 427254 138204 462698
rect 137604 427018 137786 427254
rect 138022 427018 138204 427254
rect 137604 426934 138204 427018
rect 137604 426698 137786 426934
rect 138022 426698 138204 426934
rect 137604 391254 138204 426698
rect 137604 391018 137786 391254
rect 138022 391018 138204 391254
rect 137604 390934 138204 391018
rect 137604 390698 137786 390934
rect 138022 390698 138204 390934
rect 137604 355254 138204 390698
rect 137604 355018 137786 355254
rect 138022 355018 138204 355254
rect 137604 354934 138204 355018
rect 137604 354698 137786 354934
rect 138022 354698 138204 354934
rect 137604 319254 138204 354698
rect 137604 319018 137786 319254
rect 138022 319018 138204 319254
rect 137604 318934 138204 319018
rect 137604 318698 137786 318934
rect 138022 318698 138204 318934
rect 137604 283254 138204 318698
rect 137604 283018 137786 283254
rect 138022 283018 138204 283254
rect 137604 282934 138204 283018
rect 137604 282698 137786 282934
rect 138022 282698 138204 282934
rect 137604 247254 138204 282698
rect 137604 247018 137786 247254
rect 138022 247018 138204 247254
rect 137604 246934 138204 247018
rect 137604 246698 137786 246934
rect 138022 246698 138204 246934
rect 137604 211254 138204 246698
rect 137604 211018 137786 211254
rect 138022 211018 138204 211254
rect 137604 210934 138204 211018
rect 137604 210698 137786 210934
rect 138022 210698 138204 210934
rect 137604 175254 138204 210698
rect 137604 175018 137786 175254
rect 138022 175018 138204 175254
rect 137604 174934 138204 175018
rect 137604 174698 137786 174934
rect 138022 174698 138204 174934
rect 137604 139254 138204 174698
rect 137604 139018 137786 139254
rect 138022 139018 138204 139254
rect 137604 138934 138204 139018
rect 137604 138698 137786 138934
rect 138022 138698 138204 138934
rect 137604 103254 138204 138698
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6102 119786 -5866
rect 120022 -6102 120204 -5866
rect 119604 -6186 120204 -6102
rect 119604 -6422 119786 -6186
rect 120022 -6422 120204 -6186
rect 119604 -7364 120204 -6422
rect 137604 -6786 138204 30698
rect 144804 704838 145404 705780
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 144804 542454 145404 577898
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 506454 145404 541898
rect 144804 506218 144986 506454
rect 145222 506218 145404 506454
rect 144804 506134 145404 506218
rect 144804 505898 144986 506134
rect 145222 505898 145404 506134
rect 144804 470454 145404 505898
rect 144804 470218 144986 470454
rect 145222 470218 145404 470454
rect 144804 470134 145404 470218
rect 144804 469898 144986 470134
rect 145222 469898 145404 470134
rect 144804 434454 145404 469898
rect 144804 434218 144986 434454
rect 145222 434218 145404 434454
rect 144804 434134 145404 434218
rect 144804 433898 144986 434134
rect 145222 433898 145404 434134
rect 144804 398454 145404 433898
rect 144804 398218 144986 398454
rect 145222 398218 145404 398454
rect 144804 398134 145404 398218
rect 144804 397898 144986 398134
rect 145222 397898 145404 398134
rect 144804 362454 145404 397898
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 326454 145404 361898
rect 144804 326218 144986 326454
rect 145222 326218 145404 326454
rect 144804 326134 145404 326218
rect 144804 325898 144986 326134
rect 145222 325898 145404 326134
rect 144804 290454 145404 325898
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 218454 145404 253898
rect 144804 218218 144986 218454
rect 145222 218218 145404 218454
rect 144804 218134 145404 218218
rect 144804 217898 144986 218134
rect 145222 217898 145404 218134
rect 144804 182454 145404 217898
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1844 145404 -902
rect 148404 690054 149004 706122
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 510054 149004 545498
rect 148404 509818 148586 510054
rect 148822 509818 149004 510054
rect 148404 509734 149004 509818
rect 148404 509498 148586 509734
rect 148822 509498 149004 509734
rect 148404 474054 149004 509498
rect 148404 473818 148586 474054
rect 148822 473818 149004 474054
rect 148404 473734 149004 473818
rect 148404 473498 148586 473734
rect 148822 473498 149004 473734
rect 148404 438054 149004 473498
rect 148404 437818 148586 438054
rect 148822 437818 149004 438054
rect 148404 437734 149004 437818
rect 148404 437498 148586 437734
rect 148822 437498 149004 437734
rect 148404 402054 149004 437498
rect 148404 401818 148586 402054
rect 148822 401818 149004 402054
rect 148404 401734 149004 401818
rect 148404 401498 148586 401734
rect 148822 401498 149004 401734
rect 148404 366054 149004 401498
rect 148404 365818 148586 366054
rect 148822 365818 149004 366054
rect 148404 365734 149004 365818
rect 148404 365498 148586 365734
rect 148822 365498 149004 365734
rect 148404 330054 149004 365498
rect 148404 329818 148586 330054
rect 148822 329818 149004 330054
rect 148404 329734 149004 329818
rect 148404 329498 148586 329734
rect 148822 329498 149004 329734
rect 148404 294054 149004 329498
rect 148404 293818 148586 294054
rect 148822 293818 149004 294054
rect 148404 293734 149004 293818
rect 148404 293498 148586 293734
rect 148822 293498 149004 293734
rect 148404 258054 149004 293498
rect 148404 257818 148586 258054
rect 148822 257818 149004 258054
rect 148404 257734 149004 257818
rect 148404 257498 148586 257734
rect 148822 257498 149004 257734
rect 148404 222054 149004 257498
rect 148404 221818 148586 222054
rect 148822 221818 149004 222054
rect 148404 221734 149004 221818
rect 148404 221498 148586 221734
rect 148822 221498 149004 221734
rect 148404 186054 149004 221498
rect 148404 185818 148586 186054
rect 148822 185818 149004 186054
rect 148404 185734 149004 185818
rect 148404 185498 148586 185734
rect 148822 185498 149004 185734
rect 148404 150054 149004 185498
rect 148404 149818 148586 150054
rect 148822 149818 149004 150054
rect 148404 149734 149004 149818
rect 148404 149498 148586 149734
rect 148822 149498 149004 149734
rect 148404 114054 149004 149498
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2186 149004 5498
rect 148404 -2422 148586 -2186
rect 148822 -2422 149004 -2186
rect 148404 -2506 149004 -2422
rect 148404 -2742 148586 -2506
rect 148822 -2742 149004 -2506
rect 148404 -3684 149004 -2742
rect 152004 693654 152604 707962
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 152004 549654 152604 585098
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 152004 513654 152604 549098
rect 152004 513418 152186 513654
rect 152422 513418 152604 513654
rect 152004 513334 152604 513418
rect 152004 513098 152186 513334
rect 152422 513098 152604 513334
rect 152004 477654 152604 513098
rect 152004 477418 152186 477654
rect 152422 477418 152604 477654
rect 152004 477334 152604 477418
rect 152004 477098 152186 477334
rect 152422 477098 152604 477334
rect 152004 441654 152604 477098
rect 152004 441418 152186 441654
rect 152422 441418 152604 441654
rect 152004 441334 152604 441418
rect 152004 441098 152186 441334
rect 152422 441098 152604 441334
rect 152004 405654 152604 441098
rect 152004 405418 152186 405654
rect 152422 405418 152604 405654
rect 152004 405334 152604 405418
rect 152004 405098 152186 405334
rect 152422 405098 152604 405334
rect 152004 369654 152604 405098
rect 152004 369418 152186 369654
rect 152422 369418 152604 369654
rect 152004 369334 152604 369418
rect 152004 369098 152186 369334
rect 152422 369098 152604 369334
rect 152004 333654 152604 369098
rect 152004 333418 152186 333654
rect 152422 333418 152604 333654
rect 152004 333334 152604 333418
rect 152004 333098 152186 333334
rect 152422 333098 152604 333334
rect 152004 297654 152604 333098
rect 152004 297418 152186 297654
rect 152422 297418 152604 297654
rect 152004 297334 152604 297418
rect 152004 297098 152186 297334
rect 152422 297098 152604 297334
rect 152004 261654 152604 297098
rect 152004 261418 152186 261654
rect 152422 261418 152604 261654
rect 152004 261334 152604 261418
rect 152004 261098 152186 261334
rect 152422 261098 152604 261334
rect 152004 225654 152604 261098
rect 152004 225418 152186 225654
rect 152422 225418 152604 225654
rect 152004 225334 152604 225418
rect 152004 225098 152186 225334
rect 152422 225098 152604 225334
rect 152004 189654 152604 225098
rect 152004 189418 152186 189654
rect 152422 189418 152604 189654
rect 152004 189334 152604 189418
rect 152004 189098 152186 189334
rect 152422 189098 152604 189334
rect 152004 153654 152604 189098
rect 152004 153418 152186 153654
rect 152422 153418 152604 153654
rect 152004 153334 152604 153418
rect 152004 153098 152186 153334
rect 152422 153098 152604 153334
rect 152004 117654 152604 153098
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4026 152604 9098
rect 152004 -4262 152186 -4026
rect 152422 -4262 152604 -4026
rect 152004 -4346 152604 -4262
rect 152004 -4582 152186 -4346
rect 152422 -4582 152604 -4346
rect 152004 -5524 152604 -4582
rect 155604 697254 156204 709802
rect 173604 711278 174204 711300
rect 173604 711042 173786 711278
rect 174022 711042 174204 711278
rect 173604 710958 174204 711042
rect 173604 710722 173786 710958
rect 174022 710722 174204 710958
rect 170004 709438 170604 709460
rect 170004 709202 170186 709438
rect 170422 709202 170604 709438
rect 170004 709118 170604 709202
rect 170004 708882 170186 709118
rect 170422 708882 170604 709118
rect 166404 707598 167004 707620
rect 166404 707362 166586 707598
rect 166822 707362 167004 707598
rect 166404 707278 167004 707362
rect 166404 707042 166586 707278
rect 166822 707042 167004 707278
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 155604 553254 156204 588698
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 155604 517254 156204 552698
rect 155604 517018 155786 517254
rect 156022 517018 156204 517254
rect 155604 516934 156204 517018
rect 155604 516698 155786 516934
rect 156022 516698 156204 516934
rect 155604 481254 156204 516698
rect 155604 481018 155786 481254
rect 156022 481018 156204 481254
rect 155604 480934 156204 481018
rect 155604 480698 155786 480934
rect 156022 480698 156204 480934
rect 155604 445254 156204 480698
rect 155604 445018 155786 445254
rect 156022 445018 156204 445254
rect 155604 444934 156204 445018
rect 155604 444698 155786 444934
rect 156022 444698 156204 444934
rect 155604 409254 156204 444698
rect 155604 409018 155786 409254
rect 156022 409018 156204 409254
rect 155604 408934 156204 409018
rect 155604 408698 155786 408934
rect 156022 408698 156204 408934
rect 155604 373254 156204 408698
rect 155604 373018 155786 373254
rect 156022 373018 156204 373254
rect 155604 372934 156204 373018
rect 155604 372698 155786 372934
rect 156022 372698 156204 372934
rect 155604 337254 156204 372698
rect 155604 337018 155786 337254
rect 156022 337018 156204 337254
rect 155604 336934 156204 337018
rect 155604 336698 155786 336934
rect 156022 336698 156204 336934
rect 155604 301254 156204 336698
rect 155604 301018 155786 301254
rect 156022 301018 156204 301254
rect 155604 300934 156204 301018
rect 155604 300698 155786 300934
rect 156022 300698 156204 300934
rect 155604 265254 156204 300698
rect 155604 265018 155786 265254
rect 156022 265018 156204 265254
rect 155604 264934 156204 265018
rect 155604 264698 155786 264934
rect 156022 264698 156204 264934
rect 155604 229254 156204 264698
rect 155604 229018 155786 229254
rect 156022 229018 156204 229254
rect 155604 228934 156204 229018
rect 155604 228698 155786 228934
rect 156022 228698 156204 228934
rect 155604 193254 156204 228698
rect 155604 193018 155786 193254
rect 156022 193018 156204 193254
rect 155604 192934 156204 193018
rect 155604 192698 155786 192934
rect 156022 192698 156204 192934
rect 155604 157254 156204 192698
rect 155604 157018 155786 157254
rect 156022 157018 156204 157254
rect 155604 156934 156204 157018
rect 155604 156698 155786 156934
rect 156022 156698 156204 156934
rect 155604 121254 156204 156698
rect 155604 121018 155786 121254
rect 156022 121018 156204 121254
rect 155604 120934 156204 121018
rect 155604 120698 155786 120934
rect 156022 120698 156204 120934
rect 155604 85254 156204 120698
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7022 137786 -6786
rect 138022 -7022 138204 -6786
rect 137604 -7106 138204 -7022
rect 137604 -7342 137786 -7106
rect 138022 -7342 138204 -7106
rect 137604 -7364 138204 -7342
rect 155604 -5866 156204 12698
rect 162804 705758 163404 705780
rect 162804 705522 162986 705758
rect 163222 705522 163404 705758
rect 162804 705438 163404 705522
rect 162804 705202 162986 705438
rect 163222 705202 163404 705438
rect 162804 668454 163404 705202
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 524454 163404 559898
rect 162804 524218 162986 524454
rect 163222 524218 163404 524454
rect 162804 524134 163404 524218
rect 162804 523898 162986 524134
rect 163222 523898 163404 524134
rect 162804 488454 163404 523898
rect 162804 488218 162986 488454
rect 163222 488218 163404 488454
rect 162804 488134 163404 488218
rect 162804 487898 162986 488134
rect 163222 487898 163404 488134
rect 162804 452454 163404 487898
rect 162804 452218 162986 452454
rect 163222 452218 163404 452454
rect 162804 452134 163404 452218
rect 162804 451898 162986 452134
rect 163222 451898 163404 452134
rect 162804 416454 163404 451898
rect 162804 416218 162986 416454
rect 163222 416218 163404 416454
rect 162804 416134 163404 416218
rect 162804 415898 162986 416134
rect 163222 415898 163404 416134
rect 162804 380454 163404 415898
rect 162804 380218 162986 380454
rect 163222 380218 163404 380454
rect 162804 380134 163404 380218
rect 162804 379898 162986 380134
rect 163222 379898 163404 380134
rect 162804 344454 163404 379898
rect 162804 344218 162986 344454
rect 163222 344218 163404 344454
rect 162804 344134 163404 344218
rect 162804 343898 162986 344134
rect 163222 343898 163404 344134
rect 162804 308454 163404 343898
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 272454 163404 307898
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 236454 163404 271898
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 200454 163404 235898
rect 162804 200218 162986 200454
rect 163222 200218 163404 200454
rect 162804 200134 163404 200218
rect 162804 199898 162986 200134
rect 163222 199898 163404 200134
rect 162804 164454 163404 199898
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1266 163404 19898
rect 162804 -1502 162986 -1266
rect 163222 -1502 163404 -1266
rect 162804 -1586 163404 -1502
rect 162804 -1822 162986 -1586
rect 163222 -1822 163404 -1586
rect 162804 -1844 163404 -1822
rect 166404 672054 167004 707042
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 528054 167004 563498
rect 166404 527818 166586 528054
rect 166822 527818 167004 528054
rect 166404 527734 167004 527818
rect 166404 527498 166586 527734
rect 166822 527498 167004 527734
rect 166404 492054 167004 527498
rect 166404 491818 166586 492054
rect 166822 491818 167004 492054
rect 166404 491734 167004 491818
rect 166404 491498 166586 491734
rect 166822 491498 167004 491734
rect 166404 456054 167004 491498
rect 166404 455818 166586 456054
rect 166822 455818 167004 456054
rect 166404 455734 167004 455818
rect 166404 455498 166586 455734
rect 166822 455498 167004 455734
rect 166404 420054 167004 455498
rect 166404 419818 166586 420054
rect 166822 419818 167004 420054
rect 166404 419734 167004 419818
rect 166404 419498 166586 419734
rect 166822 419498 167004 419734
rect 166404 384054 167004 419498
rect 166404 383818 166586 384054
rect 166822 383818 167004 384054
rect 166404 383734 167004 383818
rect 166404 383498 166586 383734
rect 166822 383498 167004 383734
rect 166404 348054 167004 383498
rect 166404 347818 166586 348054
rect 166822 347818 167004 348054
rect 166404 347734 167004 347818
rect 166404 347498 166586 347734
rect 166822 347498 167004 347734
rect 166404 312054 167004 347498
rect 166404 311818 166586 312054
rect 166822 311818 167004 312054
rect 166404 311734 167004 311818
rect 166404 311498 166586 311734
rect 166822 311498 167004 311734
rect 166404 276054 167004 311498
rect 166404 275818 166586 276054
rect 166822 275818 167004 276054
rect 166404 275734 167004 275818
rect 166404 275498 166586 275734
rect 166822 275498 167004 275734
rect 166404 240054 167004 275498
rect 166404 239818 166586 240054
rect 166822 239818 167004 240054
rect 166404 239734 167004 239818
rect 166404 239498 166586 239734
rect 166822 239498 167004 239734
rect 166404 204054 167004 239498
rect 166404 203818 166586 204054
rect 166822 203818 167004 204054
rect 166404 203734 167004 203818
rect 166404 203498 166586 203734
rect 166822 203498 167004 203734
rect 166404 168054 167004 203498
rect 166404 167818 166586 168054
rect 166822 167818 167004 168054
rect 166404 167734 167004 167818
rect 166404 167498 166586 167734
rect 166822 167498 167004 167734
rect 166404 132054 167004 167498
rect 166404 131818 166586 132054
rect 166822 131818 167004 132054
rect 166404 131734 167004 131818
rect 166404 131498 166586 131734
rect 166822 131498 167004 131734
rect 166404 96054 167004 131498
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3106 167004 23498
rect 166404 -3342 166586 -3106
rect 166822 -3342 167004 -3106
rect 166404 -3426 167004 -3342
rect 166404 -3662 166586 -3426
rect 166822 -3662 167004 -3426
rect 166404 -3684 167004 -3662
rect 170004 675654 170604 708882
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 170004 531654 170604 567098
rect 170004 531418 170186 531654
rect 170422 531418 170604 531654
rect 170004 531334 170604 531418
rect 170004 531098 170186 531334
rect 170422 531098 170604 531334
rect 170004 495654 170604 531098
rect 170004 495418 170186 495654
rect 170422 495418 170604 495654
rect 170004 495334 170604 495418
rect 170004 495098 170186 495334
rect 170422 495098 170604 495334
rect 170004 459654 170604 495098
rect 170004 459418 170186 459654
rect 170422 459418 170604 459654
rect 170004 459334 170604 459418
rect 170004 459098 170186 459334
rect 170422 459098 170604 459334
rect 170004 423654 170604 459098
rect 170004 423418 170186 423654
rect 170422 423418 170604 423654
rect 170004 423334 170604 423418
rect 170004 423098 170186 423334
rect 170422 423098 170604 423334
rect 170004 387654 170604 423098
rect 170004 387418 170186 387654
rect 170422 387418 170604 387654
rect 170004 387334 170604 387418
rect 170004 387098 170186 387334
rect 170422 387098 170604 387334
rect 170004 351654 170604 387098
rect 170004 351418 170186 351654
rect 170422 351418 170604 351654
rect 170004 351334 170604 351418
rect 170004 351098 170186 351334
rect 170422 351098 170604 351334
rect 170004 315654 170604 351098
rect 170004 315418 170186 315654
rect 170422 315418 170604 315654
rect 170004 315334 170604 315418
rect 170004 315098 170186 315334
rect 170422 315098 170604 315334
rect 170004 279654 170604 315098
rect 170004 279418 170186 279654
rect 170422 279418 170604 279654
rect 170004 279334 170604 279418
rect 170004 279098 170186 279334
rect 170422 279098 170604 279334
rect 170004 243654 170604 279098
rect 170004 243418 170186 243654
rect 170422 243418 170604 243654
rect 170004 243334 170604 243418
rect 170004 243098 170186 243334
rect 170422 243098 170604 243334
rect 170004 207654 170604 243098
rect 170004 207418 170186 207654
rect 170422 207418 170604 207654
rect 170004 207334 170604 207418
rect 170004 207098 170186 207334
rect 170422 207098 170604 207334
rect 170004 171654 170604 207098
rect 170004 171418 170186 171654
rect 170422 171418 170604 171654
rect 170004 171334 170604 171418
rect 170004 171098 170186 171334
rect 170422 171098 170604 171334
rect 170004 135654 170604 171098
rect 170004 135418 170186 135654
rect 170422 135418 170604 135654
rect 170004 135334 170604 135418
rect 170004 135098 170186 135334
rect 170422 135098 170604 135334
rect 170004 99654 170604 135098
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -4946 170604 27098
rect 170004 -5182 170186 -4946
rect 170422 -5182 170604 -4946
rect 170004 -5266 170604 -5182
rect 170004 -5502 170186 -5266
rect 170422 -5502 170604 -5266
rect 170004 -5524 170604 -5502
rect 173604 679254 174204 710722
rect 191604 710358 192204 711300
rect 191604 710122 191786 710358
rect 192022 710122 192204 710358
rect 191604 710038 192204 710122
rect 191604 709802 191786 710038
rect 192022 709802 192204 710038
rect 188004 708518 188604 709460
rect 188004 708282 188186 708518
rect 188422 708282 188604 708518
rect 188004 708198 188604 708282
rect 188004 707962 188186 708198
rect 188422 707962 188604 708198
rect 184404 706678 185004 707620
rect 184404 706442 184586 706678
rect 184822 706442 185004 706678
rect 184404 706358 185004 706442
rect 184404 706122 184586 706358
rect 184822 706122 185004 706358
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 535254 174204 570698
rect 173604 535018 173786 535254
rect 174022 535018 174204 535254
rect 173604 534934 174204 535018
rect 173604 534698 173786 534934
rect 174022 534698 174204 534934
rect 173604 499254 174204 534698
rect 173604 499018 173786 499254
rect 174022 499018 174204 499254
rect 173604 498934 174204 499018
rect 173604 498698 173786 498934
rect 174022 498698 174204 498934
rect 173604 463254 174204 498698
rect 173604 463018 173786 463254
rect 174022 463018 174204 463254
rect 173604 462934 174204 463018
rect 173604 462698 173786 462934
rect 174022 462698 174204 462934
rect 173604 427254 174204 462698
rect 173604 427018 173786 427254
rect 174022 427018 174204 427254
rect 173604 426934 174204 427018
rect 173604 426698 173786 426934
rect 174022 426698 174204 426934
rect 173604 391254 174204 426698
rect 173604 391018 173786 391254
rect 174022 391018 174204 391254
rect 173604 390934 174204 391018
rect 173604 390698 173786 390934
rect 174022 390698 174204 390934
rect 173604 355254 174204 390698
rect 173604 355018 173786 355254
rect 174022 355018 174204 355254
rect 173604 354934 174204 355018
rect 173604 354698 173786 354934
rect 174022 354698 174204 354934
rect 173604 319254 174204 354698
rect 173604 319018 173786 319254
rect 174022 319018 174204 319254
rect 173604 318934 174204 319018
rect 173604 318698 173786 318934
rect 174022 318698 174204 318934
rect 173604 283254 174204 318698
rect 173604 283018 173786 283254
rect 174022 283018 174204 283254
rect 173604 282934 174204 283018
rect 173604 282698 173786 282934
rect 174022 282698 174204 282934
rect 173604 247254 174204 282698
rect 173604 247018 173786 247254
rect 174022 247018 174204 247254
rect 173604 246934 174204 247018
rect 173604 246698 173786 246934
rect 174022 246698 174204 246934
rect 173604 211254 174204 246698
rect 173604 211018 173786 211254
rect 174022 211018 174204 211254
rect 173604 210934 174204 211018
rect 173604 210698 173786 210934
rect 174022 210698 174204 210934
rect 173604 175254 174204 210698
rect 173604 175018 173786 175254
rect 174022 175018 174204 175254
rect 173604 174934 174204 175018
rect 173604 174698 173786 174934
rect 174022 174698 174204 174934
rect 173604 139254 174204 174698
rect 173604 139018 173786 139254
rect 174022 139018 174204 139254
rect 173604 138934 174204 139018
rect 173604 138698 173786 138934
rect 174022 138698 174204 138934
rect 173604 103254 174204 138698
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6102 155786 -5866
rect 156022 -6102 156204 -5866
rect 155604 -6186 156204 -6102
rect 155604 -6422 155786 -6186
rect 156022 -6422 156204 -6186
rect 155604 -7364 156204 -6422
rect 173604 -6786 174204 30698
rect 180804 704838 181404 705780
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 506454 181404 541898
rect 180804 506218 180986 506454
rect 181222 506218 181404 506454
rect 180804 506134 181404 506218
rect 180804 505898 180986 506134
rect 181222 505898 181404 506134
rect 180804 470454 181404 505898
rect 180804 470218 180986 470454
rect 181222 470218 181404 470454
rect 180804 470134 181404 470218
rect 180804 469898 180986 470134
rect 181222 469898 181404 470134
rect 180804 434454 181404 469898
rect 180804 434218 180986 434454
rect 181222 434218 181404 434454
rect 180804 434134 181404 434218
rect 180804 433898 180986 434134
rect 181222 433898 181404 434134
rect 180804 398454 181404 433898
rect 180804 398218 180986 398454
rect 181222 398218 181404 398454
rect 180804 398134 181404 398218
rect 180804 397898 180986 398134
rect 181222 397898 181404 398134
rect 180804 362454 181404 397898
rect 180804 362218 180986 362454
rect 181222 362218 181404 362454
rect 180804 362134 181404 362218
rect 180804 361898 180986 362134
rect 181222 361898 181404 362134
rect 180804 326454 181404 361898
rect 180804 326218 180986 326454
rect 181222 326218 181404 326454
rect 180804 326134 181404 326218
rect 180804 325898 180986 326134
rect 181222 325898 181404 326134
rect 180804 290454 181404 325898
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 254454 181404 289898
rect 180804 254218 180986 254454
rect 181222 254218 181404 254454
rect 180804 254134 181404 254218
rect 180804 253898 180986 254134
rect 181222 253898 181404 254134
rect 180804 218454 181404 253898
rect 180804 218218 180986 218454
rect 181222 218218 181404 218454
rect 180804 218134 181404 218218
rect 180804 217898 180986 218134
rect 181222 217898 181404 218134
rect 180804 182454 181404 217898
rect 180804 182218 180986 182454
rect 181222 182218 181404 182454
rect 180804 182134 181404 182218
rect 180804 181898 180986 182134
rect 181222 181898 181404 182134
rect 180804 146454 181404 181898
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1844 181404 -902
rect 184404 690054 185004 706122
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 510054 185004 545498
rect 184404 509818 184586 510054
rect 184822 509818 185004 510054
rect 184404 509734 185004 509818
rect 184404 509498 184586 509734
rect 184822 509498 185004 509734
rect 184404 474054 185004 509498
rect 184404 473818 184586 474054
rect 184822 473818 185004 474054
rect 184404 473734 185004 473818
rect 184404 473498 184586 473734
rect 184822 473498 185004 473734
rect 184404 438054 185004 473498
rect 184404 437818 184586 438054
rect 184822 437818 185004 438054
rect 184404 437734 185004 437818
rect 184404 437498 184586 437734
rect 184822 437498 185004 437734
rect 184404 402054 185004 437498
rect 184404 401818 184586 402054
rect 184822 401818 185004 402054
rect 184404 401734 185004 401818
rect 184404 401498 184586 401734
rect 184822 401498 185004 401734
rect 184404 366054 185004 401498
rect 184404 365818 184586 366054
rect 184822 365818 185004 366054
rect 184404 365734 185004 365818
rect 184404 365498 184586 365734
rect 184822 365498 185004 365734
rect 184404 330054 185004 365498
rect 184404 329818 184586 330054
rect 184822 329818 185004 330054
rect 184404 329734 185004 329818
rect 184404 329498 184586 329734
rect 184822 329498 185004 329734
rect 184404 294054 185004 329498
rect 184404 293818 184586 294054
rect 184822 293818 185004 294054
rect 184404 293734 185004 293818
rect 184404 293498 184586 293734
rect 184822 293498 185004 293734
rect 184404 258054 185004 293498
rect 184404 257818 184586 258054
rect 184822 257818 185004 258054
rect 184404 257734 185004 257818
rect 184404 257498 184586 257734
rect 184822 257498 185004 257734
rect 184404 222054 185004 257498
rect 184404 221818 184586 222054
rect 184822 221818 185004 222054
rect 184404 221734 185004 221818
rect 184404 221498 184586 221734
rect 184822 221498 185004 221734
rect 184404 186054 185004 221498
rect 184404 185818 184586 186054
rect 184822 185818 185004 186054
rect 184404 185734 185004 185818
rect 184404 185498 184586 185734
rect 184822 185498 185004 185734
rect 184404 150054 185004 185498
rect 184404 149818 184586 150054
rect 184822 149818 185004 150054
rect 184404 149734 185004 149818
rect 184404 149498 184586 149734
rect 184822 149498 185004 149734
rect 184404 114054 185004 149498
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2186 185004 5498
rect 184404 -2422 184586 -2186
rect 184822 -2422 185004 -2186
rect 184404 -2506 185004 -2422
rect 184404 -2742 184586 -2506
rect 184822 -2742 185004 -2506
rect 184404 -3684 185004 -2742
rect 188004 693654 188604 707962
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 585654 188604 621098
rect 188004 585418 188186 585654
rect 188422 585418 188604 585654
rect 188004 585334 188604 585418
rect 188004 585098 188186 585334
rect 188422 585098 188604 585334
rect 188004 549654 188604 585098
rect 188004 549418 188186 549654
rect 188422 549418 188604 549654
rect 188004 549334 188604 549418
rect 188004 549098 188186 549334
rect 188422 549098 188604 549334
rect 188004 513654 188604 549098
rect 188004 513418 188186 513654
rect 188422 513418 188604 513654
rect 188004 513334 188604 513418
rect 188004 513098 188186 513334
rect 188422 513098 188604 513334
rect 188004 477654 188604 513098
rect 188004 477418 188186 477654
rect 188422 477418 188604 477654
rect 188004 477334 188604 477418
rect 188004 477098 188186 477334
rect 188422 477098 188604 477334
rect 188004 441654 188604 477098
rect 188004 441418 188186 441654
rect 188422 441418 188604 441654
rect 188004 441334 188604 441418
rect 188004 441098 188186 441334
rect 188422 441098 188604 441334
rect 188004 405654 188604 441098
rect 188004 405418 188186 405654
rect 188422 405418 188604 405654
rect 188004 405334 188604 405418
rect 188004 405098 188186 405334
rect 188422 405098 188604 405334
rect 188004 369654 188604 405098
rect 188004 369418 188186 369654
rect 188422 369418 188604 369654
rect 188004 369334 188604 369418
rect 188004 369098 188186 369334
rect 188422 369098 188604 369334
rect 188004 333654 188604 369098
rect 188004 333418 188186 333654
rect 188422 333418 188604 333654
rect 188004 333334 188604 333418
rect 188004 333098 188186 333334
rect 188422 333098 188604 333334
rect 188004 297654 188604 333098
rect 188004 297418 188186 297654
rect 188422 297418 188604 297654
rect 188004 297334 188604 297418
rect 188004 297098 188186 297334
rect 188422 297098 188604 297334
rect 188004 261654 188604 297098
rect 188004 261418 188186 261654
rect 188422 261418 188604 261654
rect 188004 261334 188604 261418
rect 188004 261098 188186 261334
rect 188422 261098 188604 261334
rect 188004 225654 188604 261098
rect 188004 225418 188186 225654
rect 188422 225418 188604 225654
rect 188004 225334 188604 225418
rect 188004 225098 188186 225334
rect 188422 225098 188604 225334
rect 188004 189654 188604 225098
rect 188004 189418 188186 189654
rect 188422 189418 188604 189654
rect 188004 189334 188604 189418
rect 188004 189098 188186 189334
rect 188422 189098 188604 189334
rect 188004 153654 188604 189098
rect 188004 153418 188186 153654
rect 188422 153418 188604 153654
rect 188004 153334 188604 153418
rect 188004 153098 188186 153334
rect 188422 153098 188604 153334
rect 188004 117654 188604 153098
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4026 188604 9098
rect 188004 -4262 188186 -4026
rect 188422 -4262 188604 -4026
rect 188004 -4346 188604 -4262
rect 188004 -4582 188186 -4346
rect 188422 -4582 188604 -4346
rect 188004 -5524 188604 -4582
rect 191604 697254 192204 709802
rect 209604 711278 210204 711300
rect 209604 711042 209786 711278
rect 210022 711042 210204 711278
rect 209604 710958 210204 711042
rect 209604 710722 209786 710958
rect 210022 710722 210204 710958
rect 206004 709438 206604 709460
rect 206004 709202 206186 709438
rect 206422 709202 206604 709438
rect 206004 709118 206604 709202
rect 206004 708882 206186 709118
rect 206422 708882 206604 709118
rect 202404 707598 203004 707620
rect 202404 707362 202586 707598
rect 202822 707362 203004 707598
rect 202404 707278 203004 707362
rect 202404 707042 202586 707278
rect 202822 707042 203004 707278
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 625254 192204 660698
rect 191604 625018 191786 625254
rect 192022 625018 192204 625254
rect 191604 624934 192204 625018
rect 191604 624698 191786 624934
rect 192022 624698 192204 624934
rect 191604 589254 192204 624698
rect 191604 589018 191786 589254
rect 192022 589018 192204 589254
rect 191604 588934 192204 589018
rect 191604 588698 191786 588934
rect 192022 588698 192204 588934
rect 191604 553254 192204 588698
rect 191604 553018 191786 553254
rect 192022 553018 192204 553254
rect 191604 552934 192204 553018
rect 191604 552698 191786 552934
rect 192022 552698 192204 552934
rect 191604 517254 192204 552698
rect 191604 517018 191786 517254
rect 192022 517018 192204 517254
rect 191604 516934 192204 517018
rect 191604 516698 191786 516934
rect 192022 516698 192204 516934
rect 191604 481254 192204 516698
rect 191604 481018 191786 481254
rect 192022 481018 192204 481254
rect 191604 480934 192204 481018
rect 191604 480698 191786 480934
rect 192022 480698 192204 480934
rect 191604 445254 192204 480698
rect 191604 445018 191786 445254
rect 192022 445018 192204 445254
rect 191604 444934 192204 445018
rect 191604 444698 191786 444934
rect 192022 444698 192204 444934
rect 191604 409254 192204 444698
rect 191604 409018 191786 409254
rect 192022 409018 192204 409254
rect 191604 408934 192204 409018
rect 191604 408698 191786 408934
rect 192022 408698 192204 408934
rect 191604 373254 192204 408698
rect 191604 373018 191786 373254
rect 192022 373018 192204 373254
rect 191604 372934 192204 373018
rect 191604 372698 191786 372934
rect 192022 372698 192204 372934
rect 191604 337254 192204 372698
rect 191604 337018 191786 337254
rect 192022 337018 192204 337254
rect 191604 336934 192204 337018
rect 191604 336698 191786 336934
rect 192022 336698 192204 336934
rect 191604 301254 192204 336698
rect 191604 301018 191786 301254
rect 192022 301018 192204 301254
rect 191604 300934 192204 301018
rect 191604 300698 191786 300934
rect 192022 300698 192204 300934
rect 191604 265254 192204 300698
rect 191604 265018 191786 265254
rect 192022 265018 192204 265254
rect 191604 264934 192204 265018
rect 191604 264698 191786 264934
rect 192022 264698 192204 264934
rect 191604 229254 192204 264698
rect 191604 229018 191786 229254
rect 192022 229018 192204 229254
rect 191604 228934 192204 229018
rect 191604 228698 191786 228934
rect 192022 228698 192204 228934
rect 191604 193254 192204 228698
rect 191604 193018 191786 193254
rect 192022 193018 192204 193254
rect 191604 192934 192204 193018
rect 191604 192698 191786 192934
rect 192022 192698 192204 192934
rect 191604 157254 192204 192698
rect 191604 157018 191786 157254
rect 192022 157018 192204 157254
rect 191604 156934 192204 157018
rect 191604 156698 191786 156934
rect 192022 156698 192204 156934
rect 191604 121254 192204 156698
rect 191604 121018 191786 121254
rect 192022 121018 192204 121254
rect 191604 120934 192204 121018
rect 191604 120698 191786 120934
rect 192022 120698 192204 120934
rect 191604 85254 192204 120698
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7022 173786 -6786
rect 174022 -7022 174204 -6786
rect 173604 -7106 174204 -7022
rect 173604 -7342 173786 -7106
rect 174022 -7342 174204 -7106
rect 173604 -7364 174204 -7342
rect 191604 -5866 192204 12698
rect 198804 705758 199404 705780
rect 198804 705522 198986 705758
rect 199222 705522 199404 705758
rect 198804 705438 199404 705522
rect 198804 705202 198986 705438
rect 199222 705202 199404 705438
rect 198804 668454 199404 705202
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 560454 199404 595898
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 524454 199404 559898
rect 198804 524218 198986 524454
rect 199222 524218 199404 524454
rect 198804 524134 199404 524218
rect 198804 523898 198986 524134
rect 199222 523898 199404 524134
rect 198804 488454 199404 523898
rect 198804 488218 198986 488454
rect 199222 488218 199404 488454
rect 198804 488134 199404 488218
rect 198804 487898 198986 488134
rect 199222 487898 199404 488134
rect 198804 452454 199404 487898
rect 198804 452218 198986 452454
rect 199222 452218 199404 452454
rect 198804 452134 199404 452218
rect 198804 451898 198986 452134
rect 199222 451898 199404 452134
rect 198804 416454 199404 451898
rect 198804 416218 198986 416454
rect 199222 416218 199404 416454
rect 198804 416134 199404 416218
rect 198804 415898 198986 416134
rect 199222 415898 199404 416134
rect 198804 380454 199404 415898
rect 198804 380218 198986 380454
rect 199222 380218 199404 380454
rect 198804 380134 199404 380218
rect 198804 379898 198986 380134
rect 199222 379898 199404 380134
rect 198804 344454 199404 379898
rect 198804 344218 198986 344454
rect 199222 344218 199404 344454
rect 198804 344134 199404 344218
rect 198804 343898 198986 344134
rect 199222 343898 199404 344134
rect 198804 308454 199404 343898
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 272454 199404 307898
rect 198804 272218 198986 272454
rect 199222 272218 199404 272454
rect 198804 272134 199404 272218
rect 198804 271898 198986 272134
rect 199222 271898 199404 272134
rect 198804 236454 199404 271898
rect 198804 236218 198986 236454
rect 199222 236218 199404 236454
rect 198804 236134 199404 236218
rect 198804 235898 198986 236134
rect 199222 235898 199404 236134
rect 198804 200454 199404 235898
rect 198804 200218 198986 200454
rect 199222 200218 199404 200454
rect 198804 200134 199404 200218
rect 198804 199898 198986 200134
rect 199222 199898 199404 200134
rect 198804 164454 199404 199898
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1266 199404 19898
rect 198804 -1502 198986 -1266
rect 199222 -1502 199404 -1266
rect 198804 -1586 199404 -1502
rect 198804 -1822 198986 -1586
rect 199222 -1822 199404 -1586
rect 198804 -1844 199404 -1822
rect 202404 672054 203004 707042
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 600054 203004 635498
rect 202404 599818 202586 600054
rect 202822 599818 203004 600054
rect 202404 599734 203004 599818
rect 202404 599498 202586 599734
rect 202822 599498 203004 599734
rect 202404 564054 203004 599498
rect 202404 563818 202586 564054
rect 202822 563818 203004 564054
rect 202404 563734 203004 563818
rect 202404 563498 202586 563734
rect 202822 563498 203004 563734
rect 202404 528054 203004 563498
rect 202404 527818 202586 528054
rect 202822 527818 203004 528054
rect 202404 527734 203004 527818
rect 202404 527498 202586 527734
rect 202822 527498 203004 527734
rect 202404 492054 203004 527498
rect 202404 491818 202586 492054
rect 202822 491818 203004 492054
rect 202404 491734 203004 491818
rect 202404 491498 202586 491734
rect 202822 491498 203004 491734
rect 202404 456054 203004 491498
rect 202404 455818 202586 456054
rect 202822 455818 203004 456054
rect 202404 455734 203004 455818
rect 202404 455498 202586 455734
rect 202822 455498 203004 455734
rect 202404 420054 203004 455498
rect 202404 419818 202586 420054
rect 202822 419818 203004 420054
rect 202404 419734 203004 419818
rect 202404 419498 202586 419734
rect 202822 419498 203004 419734
rect 202404 384054 203004 419498
rect 202404 383818 202586 384054
rect 202822 383818 203004 384054
rect 202404 383734 203004 383818
rect 202404 383498 202586 383734
rect 202822 383498 203004 383734
rect 202404 348054 203004 383498
rect 202404 347818 202586 348054
rect 202822 347818 203004 348054
rect 202404 347734 203004 347818
rect 202404 347498 202586 347734
rect 202822 347498 203004 347734
rect 202404 312054 203004 347498
rect 202404 311818 202586 312054
rect 202822 311818 203004 312054
rect 202404 311734 203004 311818
rect 202404 311498 202586 311734
rect 202822 311498 203004 311734
rect 202404 276054 203004 311498
rect 202404 275818 202586 276054
rect 202822 275818 203004 276054
rect 202404 275734 203004 275818
rect 202404 275498 202586 275734
rect 202822 275498 203004 275734
rect 202404 240054 203004 275498
rect 202404 239818 202586 240054
rect 202822 239818 203004 240054
rect 202404 239734 203004 239818
rect 202404 239498 202586 239734
rect 202822 239498 203004 239734
rect 202404 204054 203004 239498
rect 202404 203818 202586 204054
rect 202822 203818 203004 204054
rect 202404 203734 203004 203818
rect 202404 203498 202586 203734
rect 202822 203498 203004 203734
rect 202404 168054 203004 203498
rect 202404 167818 202586 168054
rect 202822 167818 203004 168054
rect 202404 167734 203004 167818
rect 202404 167498 202586 167734
rect 202822 167498 203004 167734
rect 202404 132054 203004 167498
rect 202404 131818 202586 132054
rect 202822 131818 203004 132054
rect 202404 131734 203004 131818
rect 202404 131498 202586 131734
rect 202822 131498 203004 131734
rect 202404 96054 203004 131498
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3106 203004 23498
rect 202404 -3342 202586 -3106
rect 202822 -3342 203004 -3106
rect 202404 -3426 203004 -3342
rect 202404 -3662 202586 -3426
rect 202822 -3662 203004 -3426
rect 202404 -3684 203004 -3662
rect 206004 675654 206604 708882
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 639654 206604 675098
rect 206004 639418 206186 639654
rect 206422 639418 206604 639654
rect 206004 639334 206604 639418
rect 206004 639098 206186 639334
rect 206422 639098 206604 639334
rect 206004 603654 206604 639098
rect 206004 603418 206186 603654
rect 206422 603418 206604 603654
rect 206004 603334 206604 603418
rect 206004 603098 206186 603334
rect 206422 603098 206604 603334
rect 206004 567654 206604 603098
rect 206004 567418 206186 567654
rect 206422 567418 206604 567654
rect 206004 567334 206604 567418
rect 206004 567098 206186 567334
rect 206422 567098 206604 567334
rect 206004 531654 206604 567098
rect 206004 531418 206186 531654
rect 206422 531418 206604 531654
rect 206004 531334 206604 531418
rect 206004 531098 206186 531334
rect 206422 531098 206604 531334
rect 206004 495654 206604 531098
rect 206004 495418 206186 495654
rect 206422 495418 206604 495654
rect 206004 495334 206604 495418
rect 206004 495098 206186 495334
rect 206422 495098 206604 495334
rect 206004 459654 206604 495098
rect 206004 459418 206186 459654
rect 206422 459418 206604 459654
rect 206004 459334 206604 459418
rect 206004 459098 206186 459334
rect 206422 459098 206604 459334
rect 206004 423654 206604 459098
rect 206004 423418 206186 423654
rect 206422 423418 206604 423654
rect 206004 423334 206604 423418
rect 206004 423098 206186 423334
rect 206422 423098 206604 423334
rect 206004 387654 206604 423098
rect 206004 387418 206186 387654
rect 206422 387418 206604 387654
rect 206004 387334 206604 387418
rect 206004 387098 206186 387334
rect 206422 387098 206604 387334
rect 206004 351654 206604 387098
rect 206004 351418 206186 351654
rect 206422 351418 206604 351654
rect 206004 351334 206604 351418
rect 206004 351098 206186 351334
rect 206422 351098 206604 351334
rect 206004 315654 206604 351098
rect 206004 315418 206186 315654
rect 206422 315418 206604 315654
rect 206004 315334 206604 315418
rect 206004 315098 206186 315334
rect 206422 315098 206604 315334
rect 206004 279654 206604 315098
rect 206004 279418 206186 279654
rect 206422 279418 206604 279654
rect 206004 279334 206604 279418
rect 206004 279098 206186 279334
rect 206422 279098 206604 279334
rect 206004 243654 206604 279098
rect 206004 243418 206186 243654
rect 206422 243418 206604 243654
rect 206004 243334 206604 243418
rect 206004 243098 206186 243334
rect 206422 243098 206604 243334
rect 206004 207654 206604 243098
rect 206004 207418 206186 207654
rect 206422 207418 206604 207654
rect 206004 207334 206604 207418
rect 206004 207098 206186 207334
rect 206422 207098 206604 207334
rect 206004 171654 206604 207098
rect 206004 171418 206186 171654
rect 206422 171418 206604 171654
rect 206004 171334 206604 171418
rect 206004 171098 206186 171334
rect 206422 171098 206604 171334
rect 206004 135654 206604 171098
rect 206004 135418 206186 135654
rect 206422 135418 206604 135654
rect 206004 135334 206604 135418
rect 206004 135098 206186 135334
rect 206422 135098 206604 135334
rect 206004 99654 206604 135098
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -4946 206604 27098
rect 206004 -5182 206186 -4946
rect 206422 -5182 206604 -4946
rect 206004 -5266 206604 -5182
rect 206004 -5502 206186 -5266
rect 206422 -5502 206604 -5266
rect 206004 -5524 206604 -5502
rect 209604 679254 210204 710722
rect 227604 710358 228204 711300
rect 227604 710122 227786 710358
rect 228022 710122 228204 710358
rect 227604 710038 228204 710122
rect 227604 709802 227786 710038
rect 228022 709802 228204 710038
rect 224004 708518 224604 709460
rect 224004 708282 224186 708518
rect 224422 708282 224604 708518
rect 224004 708198 224604 708282
rect 224004 707962 224186 708198
rect 224422 707962 224604 708198
rect 220404 706678 221004 707620
rect 220404 706442 220586 706678
rect 220822 706442 221004 706678
rect 220404 706358 221004 706442
rect 220404 706122 220586 706358
rect 220822 706122 221004 706358
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 643254 210204 678698
rect 209604 643018 209786 643254
rect 210022 643018 210204 643254
rect 209604 642934 210204 643018
rect 209604 642698 209786 642934
rect 210022 642698 210204 642934
rect 209604 607254 210204 642698
rect 209604 607018 209786 607254
rect 210022 607018 210204 607254
rect 209604 606934 210204 607018
rect 209604 606698 209786 606934
rect 210022 606698 210204 606934
rect 209604 571254 210204 606698
rect 209604 571018 209786 571254
rect 210022 571018 210204 571254
rect 209604 570934 210204 571018
rect 209604 570698 209786 570934
rect 210022 570698 210204 570934
rect 209604 535254 210204 570698
rect 209604 535018 209786 535254
rect 210022 535018 210204 535254
rect 209604 534934 210204 535018
rect 209604 534698 209786 534934
rect 210022 534698 210204 534934
rect 209604 499254 210204 534698
rect 209604 499018 209786 499254
rect 210022 499018 210204 499254
rect 209604 498934 210204 499018
rect 209604 498698 209786 498934
rect 210022 498698 210204 498934
rect 209604 463254 210204 498698
rect 209604 463018 209786 463254
rect 210022 463018 210204 463254
rect 209604 462934 210204 463018
rect 209604 462698 209786 462934
rect 210022 462698 210204 462934
rect 209604 427254 210204 462698
rect 209604 427018 209786 427254
rect 210022 427018 210204 427254
rect 209604 426934 210204 427018
rect 209604 426698 209786 426934
rect 210022 426698 210204 426934
rect 209604 391254 210204 426698
rect 209604 391018 209786 391254
rect 210022 391018 210204 391254
rect 209604 390934 210204 391018
rect 209604 390698 209786 390934
rect 210022 390698 210204 390934
rect 209604 355254 210204 390698
rect 209604 355018 209786 355254
rect 210022 355018 210204 355254
rect 209604 354934 210204 355018
rect 209604 354698 209786 354934
rect 210022 354698 210204 354934
rect 209604 319254 210204 354698
rect 209604 319018 209786 319254
rect 210022 319018 210204 319254
rect 209604 318934 210204 319018
rect 209604 318698 209786 318934
rect 210022 318698 210204 318934
rect 209604 283254 210204 318698
rect 209604 283018 209786 283254
rect 210022 283018 210204 283254
rect 209604 282934 210204 283018
rect 209604 282698 209786 282934
rect 210022 282698 210204 282934
rect 209604 247254 210204 282698
rect 209604 247018 209786 247254
rect 210022 247018 210204 247254
rect 209604 246934 210204 247018
rect 209604 246698 209786 246934
rect 210022 246698 210204 246934
rect 209604 211254 210204 246698
rect 209604 211018 209786 211254
rect 210022 211018 210204 211254
rect 209604 210934 210204 211018
rect 209604 210698 209786 210934
rect 210022 210698 210204 210934
rect 209604 175254 210204 210698
rect 209604 175018 209786 175254
rect 210022 175018 210204 175254
rect 209604 174934 210204 175018
rect 209604 174698 209786 174934
rect 210022 174698 210204 174934
rect 209604 139254 210204 174698
rect 209604 139018 209786 139254
rect 210022 139018 210204 139254
rect 209604 138934 210204 139018
rect 209604 138698 209786 138934
rect 210022 138698 210204 138934
rect 209604 103254 210204 138698
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6102 191786 -5866
rect 192022 -6102 192204 -5866
rect 191604 -6186 192204 -6102
rect 191604 -6422 191786 -6186
rect 192022 -6422 192204 -6186
rect 191604 -7364 192204 -6422
rect 209604 -6786 210204 30698
rect 216804 704838 217404 705780
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 578454 217404 613898
rect 216804 578218 216986 578454
rect 217222 578218 217404 578454
rect 216804 578134 217404 578218
rect 216804 577898 216986 578134
rect 217222 577898 217404 578134
rect 216804 542454 217404 577898
rect 216804 542218 216986 542454
rect 217222 542218 217404 542454
rect 216804 542134 217404 542218
rect 216804 541898 216986 542134
rect 217222 541898 217404 542134
rect 216804 506454 217404 541898
rect 216804 506218 216986 506454
rect 217222 506218 217404 506454
rect 216804 506134 217404 506218
rect 216804 505898 216986 506134
rect 217222 505898 217404 506134
rect 216804 470454 217404 505898
rect 216804 470218 216986 470454
rect 217222 470218 217404 470454
rect 216804 470134 217404 470218
rect 216804 469898 216986 470134
rect 217222 469898 217404 470134
rect 216804 434454 217404 469898
rect 216804 434218 216986 434454
rect 217222 434218 217404 434454
rect 216804 434134 217404 434218
rect 216804 433898 216986 434134
rect 217222 433898 217404 434134
rect 216804 398454 217404 433898
rect 216804 398218 216986 398454
rect 217222 398218 217404 398454
rect 216804 398134 217404 398218
rect 216804 397898 216986 398134
rect 217222 397898 217404 398134
rect 216804 362454 217404 397898
rect 216804 362218 216986 362454
rect 217222 362218 217404 362454
rect 216804 362134 217404 362218
rect 216804 361898 216986 362134
rect 217222 361898 217404 362134
rect 216804 326454 217404 361898
rect 216804 326218 216986 326454
rect 217222 326218 217404 326454
rect 216804 326134 217404 326218
rect 216804 325898 216986 326134
rect 217222 325898 217404 326134
rect 216804 290454 217404 325898
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 254454 217404 289898
rect 216804 254218 216986 254454
rect 217222 254218 217404 254454
rect 216804 254134 217404 254218
rect 216804 253898 216986 254134
rect 217222 253898 217404 254134
rect 216804 218454 217404 253898
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 216804 182454 217404 217898
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 216804 146454 217404 181898
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1844 217404 -902
rect 220404 690054 221004 706122
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 582054 221004 617498
rect 220404 581818 220586 582054
rect 220822 581818 221004 582054
rect 220404 581734 221004 581818
rect 220404 581498 220586 581734
rect 220822 581498 221004 581734
rect 220404 546054 221004 581498
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 220404 510054 221004 545498
rect 220404 509818 220586 510054
rect 220822 509818 221004 510054
rect 220404 509734 221004 509818
rect 220404 509498 220586 509734
rect 220822 509498 221004 509734
rect 220404 474054 221004 509498
rect 220404 473818 220586 474054
rect 220822 473818 221004 474054
rect 220404 473734 221004 473818
rect 220404 473498 220586 473734
rect 220822 473498 221004 473734
rect 220404 438054 221004 473498
rect 220404 437818 220586 438054
rect 220822 437818 221004 438054
rect 220404 437734 221004 437818
rect 220404 437498 220586 437734
rect 220822 437498 221004 437734
rect 220404 402054 221004 437498
rect 220404 401818 220586 402054
rect 220822 401818 221004 402054
rect 220404 401734 221004 401818
rect 220404 401498 220586 401734
rect 220822 401498 221004 401734
rect 220404 366054 221004 401498
rect 220404 365818 220586 366054
rect 220822 365818 221004 366054
rect 220404 365734 221004 365818
rect 220404 365498 220586 365734
rect 220822 365498 221004 365734
rect 220404 330054 221004 365498
rect 220404 329818 220586 330054
rect 220822 329818 221004 330054
rect 220404 329734 221004 329818
rect 220404 329498 220586 329734
rect 220822 329498 221004 329734
rect 220404 294054 221004 329498
rect 220404 293818 220586 294054
rect 220822 293818 221004 294054
rect 220404 293734 221004 293818
rect 220404 293498 220586 293734
rect 220822 293498 221004 293734
rect 220404 258054 221004 293498
rect 220404 257818 220586 258054
rect 220822 257818 221004 258054
rect 220404 257734 221004 257818
rect 220404 257498 220586 257734
rect 220822 257498 221004 257734
rect 220404 222054 221004 257498
rect 220404 221818 220586 222054
rect 220822 221818 221004 222054
rect 220404 221734 221004 221818
rect 220404 221498 220586 221734
rect 220822 221498 221004 221734
rect 220404 186054 221004 221498
rect 220404 185818 220586 186054
rect 220822 185818 221004 186054
rect 220404 185734 221004 185818
rect 220404 185498 220586 185734
rect 220822 185498 221004 185734
rect 220404 150054 221004 185498
rect 220404 149818 220586 150054
rect 220822 149818 221004 150054
rect 220404 149734 221004 149818
rect 220404 149498 220586 149734
rect 220822 149498 221004 149734
rect 220404 114054 221004 149498
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2186 221004 5498
rect 220404 -2422 220586 -2186
rect 220822 -2422 221004 -2186
rect 220404 -2506 221004 -2422
rect 220404 -2742 220586 -2506
rect 220822 -2742 221004 -2506
rect 220404 -3684 221004 -2742
rect 224004 693654 224604 707962
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 621654 224604 657098
rect 224004 621418 224186 621654
rect 224422 621418 224604 621654
rect 224004 621334 224604 621418
rect 224004 621098 224186 621334
rect 224422 621098 224604 621334
rect 224004 585654 224604 621098
rect 224004 585418 224186 585654
rect 224422 585418 224604 585654
rect 224004 585334 224604 585418
rect 224004 585098 224186 585334
rect 224422 585098 224604 585334
rect 224004 549654 224604 585098
rect 224004 549418 224186 549654
rect 224422 549418 224604 549654
rect 224004 549334 224604 549418
rect 224004 549098 224186 549334
rect 224422 549098 224604 549334
rect 224004 513654 224604 549098
rect 224004 513418 224186 513654
rect 224422 513418 224604 513654
rect 224004 513334 224604 513418
rect 224004 513098 224186 513334
rect 224422 513098 224604 513334
rect 224004 477654 224604 513098
rect 224004 477418 224186 477654
rect 224422 477418 224604 477654
rect 224004 477334 224604 477418
rect 224004 477098 224186 477334
rect 224422 477098 224604 477334
rect 224004 441654 224604 477098
rect 224004 441418 224186 441654
rect 224422 441418 224604 441654
rect 224004 441334 224604 441418
rect 224004 441098 224186 441334
rect 224422 441098 224604 441334
rect 224004 405654 224604 441098
rect 224004 405418 224186 405654
rect 224422 405418 224604 405654
rect 224004 405334 224604 405418
rect 224004 405098 224186 405334
rect 224422 405098 224604 405334
rect 224004 369654 224604 405098
rect 224004 369418 224186 369654
rect 224422 369418 224604 369654
rect 224004 369334 224604 369418
rect 224004 369098 224186 369334
rect 224422 369098 224604 369334
rect 224004 333654 224604 369098
rect 224004 333418 224186 333654
rect 224422 333418 224604 333654
rect 224004 333334 224604 333418
rect 224004 333098 224186 333334
rect 224422 333098 224604 333334
rect 224004 297654 224604 333098
rect 224004 297418 224186 297654
rect 224422 297418 224604 297654
rect 224004 297334 224604 297418
rect 224004 297098 224186 297334
rect 224422 297098 224604 297334
rect 224004 261654 224604 297098
rect 224004 261418 224186 261654
rect 224422 261418 224604 261654
rect 224004 261334 224604 261418
rect 224004 261098 224186 261334
rect 224422 261098 224604 261334
rect 224004 225654 224604 261098
rect 224004 225418 224186 225654
rect 224422 225418 224604 225654
rect 224004 225334 224604 225418
rect 224004 225098 224186 225334
rect 224422 225098 224604 225334
rect 224004 189654 224604 225098
rect 224004 189418 224186 189654
rect 224422 189418 224604 189654
rect 224004 189334 224604 189418
rect 224004 189098 224186 189334
rect 224422 189098 224604 189334
rect 224004 153654 224604 189098
rect 224004 153418 224186 153654
rect 224422 153418 224604 153654
rect 224004 153334 224604 153418
rect 224004 153098 224186 153334
rect 224422 153098 224604 153334
rect 224004 117654 224604 153098
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4026 224604 9098
rect 224004 -4262 224186 -4026
rect 224422 -4262 224604 -4026
rect 224004 -4346 224604 -4262
rect 224004 -4582 224186 -4346
rect 224422 -4582 224604 -4346
rect 224004 -5524 224604 -4582
rect 227604 697254 228204 709802
rect 245604 711278 246204 711300
rect 245604 711042 245786 711278
rect 246022 711042 246204 711278
rect 245604 710958 246204 711042
rect 245604 710722 245786 710958
rect 246022 710722 246204 710958
rect 242004 709438 242604 709460
rect 242004 709202 242186 709438
rect 242422 709202 242604 709438
rect 242004 709118 242604 709202
rect 242004 708882 242186 709118
rect 242422 708882 242604 709118
rect 238404 707598 239004 707620
rect 238404 707362 238586 707598
rect 238822 707362 239004 707598
rect 238404 707278 239004 707362
rect 238404 707042 238586 707278
rect 238822 707042 239004 707278
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 625254 228204 660698
rect 227604 625018 227786 625254
rect 228022 625018 228204 625254
rect 227604 624934 228204 625018
rect 227604 624698 227786 624934
rect 228022 624698 228204 624934
rect 227604 589254 228204 624698
rect 227604 589018 227786 589254
rect 228022 589018 228204 589254
rect 227604 588934 228204 589018
rect 227604 588698 227786 588934
rect 228022 588698 228204 588934
rect 227604 553254 228204 588698
rect 227604 553018 227786 553254
rect 228022 553018 228204 553254
rect 227604 552934 228204 553018
rect 227604 552698 227786 552934
rect 228022 552698 228204 552934
rect 227604 517254 228204 552698
rect 227604 517018 227786 517254
rect 228022 517018 228204 517254
rect 227604 516934 228204 517018
rect 227604 516698 227786 516934
rect 228022 516698 228204 516934
rect 227604 481254 228204 516698
rect 227604 481018 227786 481254
rect 228022 481018 228204 481254
rect 227604 480934 228204 481018
rect 227604 480698 227786 480934
rect 228022 480698 228204 480934
rect 227604 445254 228204 480698
rect 234804 705758 235404 705780
rect 234804 705522 234986 705758
rect 235222 705522 235404 705758
rect 234804 705438 235404 705522
rect 234804 705202 234986 705438
rect 235222 705202 235404 705438
rect 234804 668454 235404 705202
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 234804 560454 235404 595898
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 524454 235404 559898
rect 234804 524218 234986 524454
rect 235222 524218 235404 524454
rect 234804 524134 235404 524218
rect 234804 523898 234986 524134
rect 235222 523898 235404 524134
rect 234804 488454 235404 523898
rect 234804 488218 234986 488454
rect 235222 488218 235404 488454
rect 234804 488134 235404 488218
rect 234804 487898 234986 488134
rect 235222 487898 235404 488134
rect 232451 462908 232517 462909
rect 232451 462844 232452 462908
rect 232516 462844 232517 462908
rect 232451 462843 232517 462844
rect 231715 459644 231781 459645
rect 231715 459580 231716 459644
rect 231780 459580 231781 459644
rect 231715 459579 231781 459580
rect 227604 445018 227786 445254
rect 228022 445018 228204 445254
rect 227604 444934 228204 445018
rect 227604 444698 227786 444934
rect 228022 444698 228204 444934
rect 227604 409254 228204 444698
rect 227604 409018 227786 409254
rect 228022 409018 228204 409254
rect 227604 408934 228204 409018
rect 227604 408698 227786 408934
rect 228022 408698 228204 408934
rect 227604 373254 228204 408698
rect 227604 373018 227786 373254
rect 228022 373018 228204 373254
rect 227604 372934 228204 373018
rect 227604 372698 227786 372934
rect 228022 372698 228204 372934
rect 227604 337254 228204 372698
rect 227604 337018 227786 337254
rect 228022 337018 228204 337254
rect 227604 336934 228204 337018
rect 227604 336698 227786 336934
rect 228022 336698 228204 336934
rect 227604 301254 228204 336698
rect 227604 301018 227786 301254
rect 228022 301018 228204 301254
rect 227604 300934 228204 301018
rect 227604 300698 227786 300934
rect 228022 300698 228204 300934
rect 227604 265254 228204 300698
rect 227604 265018 227786 265254
rect 228022 265018 228204 265254
rect 227604 264934 228204 265018
rect 227604 264698 227786 264934
rect 228022 264698 228204 264934
rect 227604 229254 228204 264698
rect 227604 229018 227786 229254
rect 228022 229018 228204 229254
rect 227604 228934 228204 229018
rect 227604 228698 227786 228934
rect 228022 228698 228204 228934
rect 227604 193254 228204 228698
rect 227604 193018 227786 193254
rect 228022 193018 228204 193254
rect 227604 192934 228204 193018
rect 227604 192698 227786 192934
rect 228022 192698 228204 192934
rect 227604 157254 228204 192698
rect 227604 157018 227786 157254
rect 228022 157018 228204 157254
rect 227604 156934 228204 157018
rect 227604 156698 227786 156934
rect 228022 156698 228204 156934
rect 227604 121254 228204 156698
rect 227604 121018 227786 121254
rect 228022 121018 228204 121254
rect 227604 120934 228204 121018
rect 227604 120698 227786 120934
rect 228022 120698 228204 120934
rect 227604 85254 228204 120698
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 231718 39949 231778 459579
rect 232454 452573 232514 462843
rect 233003 459644 233069 459645
rect 233003 459580 233004 459644
rect 233068 459580 233069 459644
rect 233003 459579 233069 459580
rect 233923 459644 233989 459645
rect 233923 459580 233924 459644
rect 233988 459580 233989 459644
rect 233923 459579 233989 459580
rect 232451 452572 232517 452573
rect 232451 452508 232452 452572
rect 232516 452508 232517 452572
rect 232451 452507 232517 452508
rect 232083 220828 232149 220829
rect 232083 220764 232084 220828
rect 232148 220764 232149 220828
rect 232083 220763 232149 220764
rect 232086 211173 232146 220763
rect 232083 211172 232149 211173
rect 232083 211108 232084 211172
rect 232148 211108 232149 211172
rect 232083 211107 232149 211108
rect 231715 39948 231781 39949
rect 231715 39884 231716 39948
rect 231780 39884 231781 39948
rect 231715 39883 231781 39884
rect 233006 29205 233066 459579
rect 233739 459372 233805 459373
rect 233739 459308 233740 459372
rect 233804 459308 233805 459372
rect 233739 459307 233805 459308
rect 233742 90541 233802 459307
rect 233739 90540 233805 90541
rect 233739 90476 233740 90540
rect 233804 90476 233805 90540
rect 233739 90475 233805 90476
rect 233926 63749 233986 459579
rect 234804 452454 235404 487898
rect 234804 452218 234986 452454
rect 235222 452218 235404 452454
rect 234804 452134 235404 452218
rect 234804 451898 234986 452134
rect 235222 451898 235404 452134
rect 234804 416454 235404 451898
rect 234804 416218 234986 416454
rect 235222 416218 235404 416454
rect 234804 416134 235404 416218
rect 234804 415898 234986 416134
rect 235222 415898 235404 416134
rect 234804 380454 235404 415898
rect 234804 380218 234986 380454
rect 235222 380218 235404 380454
rect 234804 380134 235404 380218
rect 234804 379898 234986 380134
rect 235222 379898 235404 380134
rect 234804 344454 235404 379898
rect 234804 344218 234986 344454
rect 235222 344218 235404 344454
rect 234804 344134 235404 344218
rect 234804 343898 234986 344134
rect 235222 343898 235404 344134
rect 234804 308454 235404 343898
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234804 272454 235404 307898
rect 234804 272218 234986 272454
rect 235222 272218 235404 272454
rect 234804 272134 235404 272218
rect 234804 271898 234986 272134
rect 235222 271898 235404 272134
rect 234804 236454 235404 271898
rect 234804 236218 234986 236454
rect 235222 236218 235404 236454
rect 234804 236134 235404 236218
rect 234804 235898 234986 236134
rect 235222 235898 235404 236134
rect 234804 200454 235404 235898
rect 234804 200218 234986 200454
rect 235222 200218 235404 200454
rect 234804 200134 235404 200218
rect 234804 199898 234986 200134
rect 235222 199898 235404 200134
rect 234804 164454 235404 199898
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 233923 63748 233989 63749
rect 233923 63684 233924 63748
rect 233988 63684 233989 63748
rect 233923 63683 233989 63684
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 233003 29204 233069 29205
rect 233003 29140 233004 29204
rect 233068 29140 233069 29204
rect 233003 29139 233069 29140
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7022 209786 -6786
rect 210022 -7022 210204 -6786
rect 209604 -7106 210204 -7022
rect 209604 -7342 209786 -7106
rect 210022 -7342 210204 -7106
rect 209604 -7364 210204 -7342
rect 227604 -5866 228204 12698
rect 234804 20454 235404 55898
rect 238404 672054 239004 707042
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 636054 239004 671498
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 600054 239004 635498
rect 238404 599818 238586 600054
rect 238822 599818 239004 600054
rect 238404 599734 239004 599818
rect 238404 599498 238586 599734
rect 238822 599498 239004 599734
rect 238404 564054 239004 599498
rect 238404 563818 238586 564054
rect 238822 563818 239004 564054
rect 238404 563734 239004 563818
rect 238404 563498 238586 563734
rect 238822 563498 239004 563734
rect 238404 528054 239004 563498
rect 238404 527818 238586 528054
rect 238822 527818 239004 528054
rect 238404 527734 239004 527818
rect 238404 527498 238586 527734
rect 238822 527498 239004 527734
rect 238404 492054 239004 527498
rect 238404 491818 238586 492054
rect 238822 491818 239004 492054
rect 238404 491734 239004 491818
rect 238404 491498 238586 491734
rect 238822 491498 239004 491734
rect 238404 456054 239004 491498
rect 238404 455818 238586 456054
rect 238822 455818 239004 456054
rect 238404 455734 239004 455818
rect 238404 455498 238586 455734
rect 238822 455498 239004 455734
rect 238404 420054 239004 455498
rect 238404 419818 238586 420054
rect 238822 419818 239004 420054
rect 238404 419734 239004 419818
rect 238404 419498 238586 419734
rect 238822 419498 239004 419734
rect 238404 384054 239004 419498
rect 238404 383818 238586 384054
rect 238822 383818 239004 384054
rect 238404 383734 239004 383818
rect 238404 383498 238586 383734
rect 238822 383498 239004 383734
rect 238404 348054 239004 383498
rect 238404 347818 238586 348054
rect 238822 347818 239004 348054
rect 238404 347734 239004 347818
rect 238404 347498 238586 347734
rect 238822 347498 239004 347734
rect 238404 312054 239004 347498
rect 238404 311818 238586 312054
rect 238822 311818 239004 312054
rect 238404 311734 239004 311818
rect 238404 311498 238586 311734
rect 238822 311498 239004 311734
rect 238404 276054 239004 311498
rect 238404 275818 238586 276054
rect 238822 275818 239004 276054
rect 238404 275734 239004 275818
rect 238404 275498 238586 275734
rect 238822 275498 239004 275734
rect 238404 240054 239004 275498
rect 238404 239818 238586 240054
rect 238822 239818 239004 240054
rect 238404 239734 239004 239818
rect 238404 239498 238586 239734
rect 238822 239498 239004 239734
rect 238404 204054 239004 239498
rect 238404 203818 238586 204054
rect 238822 203818 239004 204054
rect 238404 203734 239004 203818
rect 238404 203498 238586 203734
rect 238822 203498 239004 203734
rect 238404 168054 239004 203498
rect 238404 167818 238586 168054
rect 238822 167818 239004 168054
rect 238404 167734 239004 167818
rect 238404 167498 238586 167734
rect 238822 167498 239004 167734
rect 238404 132054 239004 167498
rect 238404 131818 238586 132054
rect 238822 131818 239004 132054
rect 238404 131734 239004 131818
rect 238404 131498 238586 131734
rect 238822 131498 239004 131734
rect 238404 96054 239004 131498
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 237419 40492 237485 40493
rect 237419 40428 237420 40492
rect 237484 40428 237485 40492
rect 237419 40427 237485 40428
rect 237422 39949 237482 40427
rect 237419 39948 237485 39949
rect 237419 39884 237420 39948
rect 237484 39884 237485 39948
rect 237419 39883 237485 39884
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1266 235404 19898
rect 234804 -1502 234986 -1266
rect 235222 -1502 235404 -1266
rect 234804 -1586 235404 -1502
rect 234804 -1822 234986 -1586
rect 235222 -1822 235404 -1586
rect 234804 -1844 235404 -1822
rect 238404 24054 239004 59498
rect 242004 675654 242604 708882
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 639654 242604 675098
rect 242004 639418 242186 639654
rect 242422 639418 242604 639654
rect 242004 639334 242604 639418
rect 242004 639098 242186 639334
rect 242422 639098 242604 639334
rect 242004 603654 242604 639098
rect 242004 603418 242186 603654
rect 242422 603418 242604 603654
rect 242004 603334 242604 603418
rect 242004 603098 242186 603334
rect 242422 603098 242604 603334
rect 242004 567654 242604 603098
rect 242004 567418 242186 567654
rect 242422 567418 242604 567654
rect 242004 567334 242604 567418
rect 242004 567098 242186 567334
rect 242422 567098 242604 567334
rect 242004 531654 242604 567098
rect 242004 531418 242186 531654
rect 242422 531418 242604 531654
rect 242004 531334 242604 531418
rect 242004 531098 242186 531334
rect 242422 531098 242604 531334
rect 242004 495654 242604 531098
rect 242004 495418 242186 495654
rect 242422 495418 242604 495654
rect 242004 495334 242604 495418
rect 242004 495098 242186 495334
rect 242422 495098 242604 495334
rect 242004 459654 242604 495098
rect 242004 459418 242186 459654
rect 242422 459418 242604 459654
rect 242004 459334 242604 459418
rect 242004 459098 242186 459334
rect 242422 459098 242604 459334
rect 242004 423654 242604 459098
rect 242004 423418 242186 423654
rect 242422 423418 242604 423654
rect 242004 423334 242604 423418
rect 242004 423098 242186 423334
rect 242422 423098 242604 423334
rect 242004 387654 242604 423098
rect 242004 387418 242186 387654
rect 242422 387418 242604 387654
rect 242004 387334 242604 387418
rect 242004 387098 242186 387334
rect 242422 387098 242604 387334
rect 242004 351654 242604 387098
rect 242004 351418 242186 351654
rect 242422 351418 242604 351654
rect 242004 351334 242604 351418
rect 242004 351098 242186 351334
rect 242422 351098 242604 351334
rect 242004 315654 242604 351098
rect 242004 315418 242186 315654
rect 242422 315418 242604 315654
rect 242004 315334 242604 315418
rect 242004 315098 242186 315334
rect 242422 315098 242604 315334
rect 242004 279654 242604 315098
rect 242004 279418 242186 279654
rect 242422 279418 242604 279654
rect 242004 279334 242604 279418
rect 242004 279098 242186 279334
rect 242422 279098 242604 279334
rect 242004 243654 242604 279098
rect 242004 243418 242186 243654
rect 242422 243418 242604 243654
rect 242004 243334 242604 243418
rect 242004 243098 242186 243334
rect 242422 243098 242604 243334
rect 242004 207654 242604 243098
rect 242004 207418 242186 207654
rect 242422 207418 242604 207654
rect 242004 207334 242604 207418
rect 242004 207098 242186 207334
rect 242422 207098 242604 207334
rect 242004 171654 242604 207098
rect 242004 171418 242186 171654
rect 242422 171418 242604 171654
rect 242004 171334 242604 171418
rect 242004 171098 242186 171334
rect 242422 171098 242604 171334
rect 242004 135654 242604 171098
rect 245604 679254 246204 710722
rect 263604 710358 264204 711300
rect 263604 710122 263786 710358
rect 264022 710122 264204 710358
rect 263604 710038 264204 710122
rect 263604 709802 263786 710038
rect 264022 709802 264204 710038
rect 260004 708518 260604 709460
rect 260004 708282 260186 708518
rect 260422 708282 260604 708518
rect 260004 708198 260604 708282
rect 260004 707962 260186 708198
rect 260422 707962 260604 708198
rect 256404 706678 257004 707620
rect 256404 706442 256586 706678
rect 256822 706442 257004 706678
rect 256404 706358 257004 706442
rect 256404 706122 256586 706358
rect 256822 706122 257004 706358
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 643254 246204 678698
rect 245604 643018 245786 643254
rect 246022 643018 246204 643254
rect 245604 642934 246204 643018
rect 245604 642698 245786 642934
rect 246022 642698 246204 642934
rect 245604 607254 246204 642698
rect 245604 607018 245786 607254
rect 246022 607018 246204 607254
rect 245604 606934 246204 607018
rect 245604 606698 245786 606934
rect 246022 606698 246204 606934
rect 245604 571254 246204 606698
rect 245604 571018 245786 571254
rect 246022 571018 246204 571254
rect 245604 570934 246204 571018
rect 245604 570698 245786 570934
rect 246022 570698 246204 570934
rect 245604 535254 246204 570698
rect 245604 535018 245786 535254
rect 246022 535018 246204 535254
rect 245604 534934 246204 535018
rect 245604 534698 245786 534934
rect 246022 534698 246204 534934
rect 245604 499254 246204 534698
rect 245604 499018 245786 499254
rect 246022 499018 246204 499254
rect 245604 498934 246204 499018
rect 245604 498698 245786 498934
rect 246022 498698 246204 498934
rect 245604 463254 246204 498698
rect 245604 463018 245786 463254
rect 246022 463018 246204 463254
rect 245604 462934 246204 463018
rect 245604 462698 245786 462934
rect 246022 462698 246204 462934
rect 245604 427254 246204 462698
rect 245604 427018 245786 427254
rect 246022 427018 246204 427254
rect 245604 426934 246204 427018
rect 245604 426698 245786 426934
rect 246022 426698 246204 426934
rect 245604 391254 246204 426698
rect 245604 391018 245786 391254
rect 246022 391018 246204 391254
rect 245604 390934 246204 391018
rect 245604 390698 245786 390934
rect 246022 390698 246204 390934
rect 245604 355254 246204 390698
rect 245604 355018 245786 355254
rect 246022 355018 246204 355254
rect 245604 354934 246204 355018
rect 245604 354698 245786 354934
rect 246022 354698 246204 354934
rect 245604 319254 246204 354698
rect 245604 319018 245786 319254
rect 246022 319018 246204 319254
rect 245604 318934 246204 319018
rect 245604 318698 245786 318934
rect 246022 318698 246204 318934
rect 245604 283254 246204 318698
rect 245604 283018 245786 283254
rect 246022 283018 246204 283254
rect 245604 282934 246204 283018
rect 245604 282698 245786 282934
rect 246022 282698 246204 282934
rect 245604 247254 246204 282698
rect 245604 247018 245786 247254
rect 246022 247018 246204 247254
rect 245604 246934 246204 247018
rect 245604 246698 245786 246934
rect 246022 246698 246204 246934
rect 245604 211254 246204 246698
rect 245604 211018 245786 211254
rect 246022 211018 246204 211254
rect 245604 210934 246204 211018
rect 245604 210698 245786 210934
rect 246022 210698 246204 210934
rect 245604 175254 246204 210698
rect 245604 175018 245786 175254
rect 246022 175018 246204 175254
rect 245604 174934 246204 175018
rect 245604 174698 245786 174934
rect 246022 174698 246204 174934
rect 245604 139254 246204 174698
rect 245604 139018 245786 139254
rect 246022 139018 246204 139254
rect 245604 138934 246204 139018
rect 245604 138698 245786 138934
rect 246022 138698 246204 138934
rect 244411 138684 244477 138685
rect 244411 138620 244412 138684
rect 244476 138620 244477 138684
rect 244411 138619 244477 138620
rect 242004 135418 242186 135654
rect 242422 135418 242604 135654
rect 242004 135334 242604 135418
rect 242004 135098 242186 135334
rect 242422 135098 242604 135334
rect 242004 99654 242604 135098
rect 244414 125629 244474 138619
rect 244411 125628 244477 125629
rect 244411 125564 244412 125628
rect 244476 125564 244477 125628
rect 244411 125563 244477 125564
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 241467 29476 241533 29477
rect 241467 29412 241468 29476
rect 241532 29412 241533 29476
rect 241467 29411 241533 29412
rect 241470 29205 241530 29411
rect 241467 29204 241533 29205
rect 241467 29140 241468 29204
rect 241532 29140 241533 29204
rect 241467 29139 241533 29140
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3106 239004 23498
rect 238404 -3342 238586 -3106
rect 238822 -3342 239004 -3106
rect 238404 -3426 239004 -3342
rect 238404 -3662 238586 -3426
rect 238822 -3662 239004 -3426
rect 238404 -3684 239004 -3662
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -4946 242604 27098
rect 242004 -5182 242186 -4946
rect 242422 -5182 242604 -4946
rect 242004 -5266 242604 -5182
rect 242004 -5502 242186 -5266
rect 242422 -5502 242604 -5266
rect 242004 -5524 242604 -5502
rect 245604 103254 246204 138698
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 245604 67254 246204 102698
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6102 227786 -5866
rect 228022 -6102 228204 -5866
rect 227604 -6186 228204 -6102
rect 227604 -6422 227786 -6186
rect 228022 -6422 228204 -6186
rect 227604 -7364 228204 -6422
rect 245604 -6786 246204 30698
rect 252804 704838 253404 705780
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 578454 253404 613898
rect 252804 578218 252986 578454
rect 253222 578218 253404 578454
rect 252804 578134 253404 578218
rect 252804 577898 252986 578134
rect 253222 577898 253404 578134
rect 252804 542454 253404 577898
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 252804 506454 253404 541898
rect 252804 506218 252986 506454
rect 253222 506218 253404 506454
rect 252804 506134 253404 506218
rect 252804 505898 252986 506134
rect 253222 505898 253404 506134
rect 252804 470454 253404 505898
rect 252804 470218 252986 470454
rect 253222 470218 253404 470454
rect 252804 470134 253404 470218
rect 252804 469898 252986 470134
rect 253222 469898 253404 470134
rect 252804 434454 253404 469898
rect 252804 434218 252986 434454
rect 253222 434218 253404 434454
rect 252804 434134 253404 434218
rect 252804 433898 252986 434134
rect 253222 433898 253404 434134
rect 252804 398454 253404 433898
rect 252804 398218 252986 398454
rect 253222 398218 253404 398454
rect 252804 398134 253404 398218
rect 252804 397898 252986 398134
rect 253222 397898 253404 398134
rect 252804 362454 253404 397898
rect 252804 362218 252986 362454
rect 253222 362218 253404 362454
rect 252804 362134 253404 362218
rect 252804 361898 252986 362134
rect 253222 361898 253404 362134
rect 252804 326454 253404 361898
rect 252804 326218 252986 326454
rect 253222 326218 253404 326454
rect 252804 326134 253404 326218
rect 252804 325898 252986 326134
rect 253222 325898 253404 326134
rect 252804 290454 253404 325898
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 252804 254454 253404 289898
rect 252804 254218 252986 254454
rect 253222 254218 253404 254454
rect 252804 254134 253404 254218
rect 252804 253898 252986 254134
rect 253222 253898 253404 254134
rect 252804 218454 253404 253898
rect 252804 218218 252986 218454
rect 253222 218218 253404 218454
rect 252804 218134 253404 218218
rect 252804 217898 252986 218134
rect 253222 217898 253404 218134
rect 252804 182454 253404 217898
rect 252804 182218 252986 182454
rect 253222 182218 253404 182454
rect 252804 182134 253404 182218
rect 252804 181898 252986 182134
rect 253222 181898 253404 182134
rect 252804 146454 253404 181898
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 252804 110454 253404 145898
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1844 253404 -902
rect 256404 690054 257004 706122
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 618054 257004 653498
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 582054 257004 617498
rect 256404 581818 256586 582054
rect 256822 581818 257004 582054
rect 256404 581734 257004 581818
rect 256404 581498 256586 581734
rect 256822 581498 257004 581734
rect 256404 546054 257004 581498
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 256404 510054 257004 545498
rect 256404 509818 256586 510054
rect 256822 509818 257004 510054
rect 256404 509734 257004 509818
rect 256404 509498 256586 509734
rect 256822 509498 257004 509734
rect 256404 474054 257004 509498
rect 256404 473818 256586 474054
rect 256822 473818 257004 474054
rect 256404 473734 257004 473818
rect 256404 473498 256586 473734
rect 256822 473498 257004 473734
rect 256404 438054 257004 473498
rect 260004 693654 260604 707962
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 621654 260604 657098
rect 260004 621418 260186 621654
rect 260422 621418 260604 621654
rect 260004 621334 260604 621418
rect 260004 621098 260186 621334
rect 260422 621098 260604 621334
rect 260004 585654 260604 621098
rect 260004 585418 260186 585654
rect 260422 585418 260604 585654
rect 260004 585334 260604 585418
rect 260004 585098 260186 585334
rect 260422 585098 260604 585334
rect 260004 549654 260604 585098
rect 260004 549418 260186 549654
rect 260422 549418 260604 549654
rect 260004 549334 260604 549418
rect 260004 549098 260186 549334
rect 260422 549098 260604 549334
rect 260004 513654 260604 549098
rect 260004 513418 260186 513654
rect 260422 513418 260604 513654
rect 260004 513334 260604 513418
rect 260004 513098 260186 513334
rect 260422 513098 260604 513334
rect 260004 477654 260604 513098
rect 260004 477418 260186 477654
rect 260422 477418 260604 477654
rect 260004 477334 260604 477418
rect 260004 477098 260186 477334
rect 260422 477098 260604 477334
rect 258947 459372 259013 459373
rect 258947 459308 258948 459372
rect 259012 459308 259013 459372
rect 258947 459307 259013 459308
rect 258950 457877 259010 459307
rect 258947 457876 259013 457877
rect 258947 457812 258948 457876
rect 259012 457812 259013 457876
rect 258947 457811 259013 457812
rect 256404 437818 256586 438054
rect 256822 437818 257004 438054
rect 256404 437734 257004 437818
rect 256404 437498 256586 437734
rect 256822 437498 257004 437734
rect 256404 402054 257004 437498
rect 256404 401818 256586 402054
rect 256822 401818 257004 402054
rect 256404 401734 257004 401818
rect 256404 401498 256586 401734
rect 256822 401498 257004 401734
rect 256404 366054 257004 401498
rect 256404 365818 256586 366054
rect 256822 365818 257004 366054
rect 256404 365734 257004 365818
rect 256404 365498 256586 365734
rect 256822 365498 257004 365734
rect 256404 330054 257004 365498
rect 256404 329818 256586 330054
rect 256822 329818 257004 330054
rect 256404 329734 257004 329818
rect 256404 329498 256586 329734
rect 256822 329498 257004 329734
rect 256404 294054 257004 329498
rect 256404 293818 256586 294054
rect 256822 293818 257004 294054
rect 256404 293734 257004 293818
rect 256404 293498 256586 293734
rect 256822 293498 257004 293734
rect 256404 258054 257004 293498
rect 256404 257818 256586 258054
rect 256822 257818 257004 258054
rect 256404 257734 257004 257818
rect 256404 257498 256586 257734
rect 256822 257498 257004 257734
rect 256404 222054 257004 257498
rect 256404 221818 256586 222054
rect 256822 221818 257004 222054
rect 256404 221734 257004 221818
rect 256404 221498 256586 221734
rect 256822 221498 257004 221734
rect 256404 186054 257004 221498
rect 256404 185818 256586 186054
rect 256822 185818 257004 186054
rect 256404 185734 257004 185818
rect 256404 185498 256586 185734
rect 256822 185498 257004 185734
rect 256404 150054 257004 185498
rect 256404 149818 256586 150054
rect 256822 149818 257004 150054
rect 256404 149734 257004 149818
rect 256404 149498 256586 149734
rect 256822 149498 257004 149734
rect 256404 114054 257004 149498
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 260004 441654 260604 477098
rect 260004 441418 260186 441654
rect 260422 441418 260604 441654
rect 260004 441334 260604 441418
rect 260004 441098 260186 441334
rect 260422 441098 260604 441334
rect 260004 405654 260604 441098
rect 260004 405418 260186 405654
rect 260422 405418 260604 405654
rect 260004 405334 260604 405418
rect 260004 405098 260186 405334
rect 260422 405098 260604 405334
rect 260004 369654 260604 405098
rect 260004 369418 260186 369654
rect 260422 369418 260604 369654
rect 260004 369334 260604 369418
rect 260004 369098 260186 369334
rect 260422 369098 260604 369334
rect 260004 333654 260604 369098
rect 260004 333418 260186 333654
rect 260422 333418 260604 333654
rect 260004 333334 260604 333418
rect 260004 333098 260186 333334
rect 260422 333098 260604 333334
rect 260004 297654 260604 333098
rect 260004 297418 260186 297654
rect 260422 297418 260604 297654
rect 260004 297334 260604 297418
rect 260004 297098 260186 297334
rect 260422 297098 260604 297334
rect 260004 261654 260604 297098
rect 260004 261418 260186 261654
rect 260422 261418 260604 261654
rect 260004 261334 260604 261418
rect 260004 261098 260186 261334
rect 260422 261098 260604 261334
rect 260004 225654 260604 261098
rect 260004 225418 260186 225654
rect 260422 225418 260604 225654
rect 260004 225334 260604 225418
rect 260004 225098 260186 225334
rect 260422 225098 260604 225334
rect 260004 189654 260604 225098
rect 260004 189418 260186 189654
rect 260422 189418 260604 189654
rect 260004 189334 260604 189418
rect 260004 189098 260186 189334
rect 260422 189098 260604 189334
rect 260004 153654 260604 189098
rect 260004 153418 260186 153654
rect 260422 153418 260604 153654
rect 260004 153334 260604 153418
rect 260004 153098 260186 153334
rect 260422 153098 260604 153334
rect 260004 117654 260604 153098
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 258027 63748 258093 63749
rect 258027 63684 258028 63748
rect 258092 63684 258093 63748
rect 258027 63683 258093 63684
rect 258030 63477 258090 63683
rect 258027 63476 258093 63477
rect 258027 63412 258028 63476
rect 258092 63412 258093 63476
rect 258027 63411 258093 63412
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2186 257004 5498
rect 256404 -2422 256586 -2186
rect 256822 -2422 257004 -2186
rect 256404 -2506 257004 -2422
rect 256404 -2742 256586 -2506
rect 256822 -2742 257004 -2506
rect 256404 -3684 257004 -2742
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4026 260604 9098
rect 260004 -4262 260186 -4026
rect 260422 -4262 260604 -4026
rect 260004 -4346 260604 -4262
rect 260004 -4582 260186 -4346
rect 260422 -4582 260604 -4346
rect 260004 -5524 260604 -4582
rect 263604 697254 264204 709802
rect 281604 711278 282204 711300
rect 281604 711042 281786 711278
rect 282022 711042 282204 711278
rect 281604 710958 282204 711042
rect 281604 710722 281786 710958
rect 282022 710722 282204 710958
rect 278004 709438 278604 709460
rect 278004 709202 278186 709438
rect 278422 709202 278604 709438
rect 278004 709118 278604 709202
rect 278004 708882 278186 709118
rect 278422 708882 278604 709118
rect 274404 707598 275004 707620
rect 274404 707362 274586 707598
rect 274822 707362 275004 707598
rect 274404 707278 275004 707362
rect 274404 707042 274586 707278
rect 274822 707042 275004 707278
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 625254 264204 660698
rect 263604 625018 263786 625254
rect 264022 625018 264204 625254
rect 263604 624934 264204 625018
rect 263604 624698 263786 624934
rect 264022 624698 264204 624934
rect 263604 589254 264204 624698
rect 263604 589018 263786 589254
rect 264022 589018 264204 589254
rect 263604 588934 264204 589018
rect 263604 588698 263786 588934
rect 264022 588698 264204 588934
rect 263604 553254 264204 588698
rect 263604 553018 263786 553254
rect 264022 553018 264204 553254
rect 263604 552934 264204 553018
rect 263604 552698 263786 552934
rect 264022 552698 264204 552934
rect 263604 517254 264204 552698
rect 263604 517018 263786 517254
rect 264022 517018 264204 517254
rect 263604 516934 264204 517018
rect 263604 516698 263786 516934
rect 264022 516698 264204 516934
rect 263604 481254 264204 516698
rect 263604 481018 263786 481254
rect 264022 481018 264204 481254
rect 263604 480934 264204 481018
rect 263604 480698 263786 480934
rect 264022 480698 264204 480934
rect 263604 445254 264204 480698
rect 263604 445018 263786 445254
rect 264022 445018 264204 445254
rect 263604 444934 264204 445018
rect 263604 444698 263786 444934
rect 264022 444698 264204 444934
rect 263604 409254 264204 444698
rect 263604 409018 263786 409254
rect 264022 409018 264204 409254
rect 263604 408934 264204 409018
rect 263604 408698 263786 408934
rect 264022 408698 264204 408934
rect 263604 373254 264204 408698
rect 263604 373018 263786 373254
rect 264022 373018 264204 373254
rect 263604 372934 264204 373018
rect 263604 372698 263786 372934
rect 264022 372698 264204 372934
rect 263604 337254 264204 372698
rect 270804 705758 271404 705780
rect 270804 705522 270986 705758
rect 271222 705522 271404 705758
rect 270804 705438 271404 705522
rect 270804 705202 270986 705438
rect 271222 705202 271404 705438
rect 270804 668454 271404 705202
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 270804 488454 271404 523898
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 270804 452454 271404 487898
rect 270804 452218 270986 452454
rect 271222 452218 271404 452454
rect 270804 452134 271404 452218
rect 270804 451898 270986 452134
rect 271222 451898 271404 452134
rect 270804 416454 271404 451898
rect 270804 416218 270986 416454
rect 271222 416218 271404 416454
rect 270804 416134 271404 416218
rect 270804 415898 270986 416134
rect 271222 415898 271404 416134
rect 270804 380454 271404 415898
rect 270804 380218 270986 380454
rect 271222 380218 271404 380454
rect 270804 380134 271404 380218
rect 270804 379898 270986 380134
rect 271222 379898 271404 380134
rect 270804 344454 271404 379898
rect 270804 344218 270986 344454
rect 271222 344218 271404 344454
rect 270804 344134 271404 344218
rect 270804 343898 270986 344134
rect 271222 343898 271404 344134
rect 266491 338060 266557 338061
rect 266491 337996 266492 338060
rect 266556 337996 266557 338060
rect 266491 337995 266557 337996
rect 263604 337018 263786 337254
rect 264022 337018 264204 337254
rect 263604 336934 264204 337018
rect 263604 336698 263786 336934
rect 264022 336698 264204 336934
rect 263604 301254 264204 336698
rect 266494 328541 266554 337995
rect 266491 328540 266557 328541
rect 266491 328476 266492 328540
rect 266556 328476 266557 328540
rect 266491 328475 266557 328476
rect 263604 301018 263786 301254
rect 264022 301018 264204 301254
rect 263604 300934 264204 301018
rect 263604 300698 263786 300934
rect 264022 300698 264204 300934
rect 263604 265254 264204 300698
rect 263604 265018 263786 265254
rect 264022 265018 264204 265254
rect 263604 264934 264204 265018
rect 263604 264698 263786 264934
rect 264022 264698 264204 264934
rect 263604 229254 264204 264698
rect 263604 229018 263786 229254
rect 264022 229018 264204 229254
rect 263604 228934 264204 229018
rect 263604 228698 263786 228934
rect 264022 228698 264204 228934
rect 263604 193254 264204 228698
rect 263604 193018 263786 193254
rect 264022 193018 264204 193254
rect 263604 192934 264204 193018
rect 263604 192698 263786 192934
rect 264022 192698 264204 192934
rect 263604 157254 264204 192698
rect 263604 157018 263786 157254
rect 264022 157018 264204 157254
rect 263604 156934 264204 157018
rect 263604 156698 263786 156934
rect 264022 156698 264204 156934
rect 263604 121254 264204 156698
rect 263604 121018 263786 121254
rect 264022 121018 264204 121254
rect 263604 120934 264204 121018
rect 263604 120698 263786 120934
rect 264022 120698 264204 120934
rect 263604 85254 264204 120698
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 270804 308454 271404 343898
rect 270804 308218 270986 308454
rect 271222 308218 271404 308454
rect 270804 308134 271404 308218
rect 270804 307898 270986 308134
rect 271222 307898 271404 308134
rect 270804 272454 271404 307898
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 270804 236454 271404 271898
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 270804 200454 271404 235898
rect 270804 200218 270986 200454
rect 271222 200218 271404 200454
rect 270804 200134 271404 200218
rect 270804 199898 270986 200134
rect 271222 199898 271404 200134
rect 270804 164454 271404 199898
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 268699 17100 268765 17101
rect 268699 17036 268700 17100
rect 268764 17036 268765 17100
rect 268699 17035 268765 17036
rect 268702 16690 268762 17035
rect 268883 16692 268949 16693
rect 268883 16690 268884 16692
rect 268702 16630 268884 16690
rect 268883 16628 268884 16630
rect 268948 16628 268949 16692
rect 268883 16627 268949 16628
rect 268883 16284 268949 16285
rect 268883 16220 268884 16284
rect 268948 16220 268949 16284
rect 268883 16219 268949 16220
rect 268886 15605 268946 16219
rect 268883 15604 268949 15605
rect 268883 15540 268884 15604
rect 268948 15540 268949 15604
rect 268883 15539 268949 15540
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7022 245786 -6786
rect 246022 -7022 246204 -6786
rect 245604 -7106 246204 -7022
rect 245604 -7342 245786 -7106
rect 246022 -7342 246204 -7106
rect 245604 -7364 246204 -7342
rect 263604 -5866 264204 12698
rect 270804 -1266 271404 19898
rect 270804 -1502 270986 -1266
rect 271222 -1502 271404 -1266
rect 270804 -1586 271404 -1502
rect 270804 -1822 270986 -1586
rect 271222 -1822 271404 -1586
rect 270804 -1844 271404 -1822
rect 274404 672054 275004 707042
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 528054 275004 563498
rect 274404 527818 274586 528054
rect 274822 527818 275004 528054
rect 274404 527734 275004 527818
rect 274404 527498 274586 527734
rect 274822 527498 275004 527734
rect 274404 492054 275004 527498
rect 274404 491818 274586 492054
rect 274822 491818 275004 492054
rect 274404 491734 275004 491818
rect 274404 491498 274586 491734
rect 274822 491498 275004 491734
rect 274404 456054 275004 491498
rect 274404 455818 274586 456054
rect 274822 455818 275004 456054
rect 274404 455734 275004 455818
rect 274404 455498 274586 455734
rect 274822 455498 275004 455734
rect 274404 420054 275004 455498
rect 274404 419818 274586 420054
rect 274822 419818 275004 420054
rect 274404 419734 275004 419818
rect 274404 419498 274586 419734
rect 274822 419498 275004 419734
rect 274404 384054 275004 419498
rect 274404 383818 274586 384054
rect 274822 383818 275004 384054
rect 274404 383734 275004 383818
rect 274404 383498 274586 383734
rect 274822 383498 275004 383734
rect 274404 348054 275004 383498
rect 274404 347818 274586 348054
rect 274822 347818 275004 348054
rect 274404 347734 275004 347818
rect 274404 347498 274586 347734
rect 274822 347498 275004 347734
rect 274404 312054 275004 347498
rect 274404 311818 274586 312054
rect 274822 311818 275004 312054
rect 274404 311734 275004 311818
rect 274404 311498 274586 311734
rect 274822 311498 275004 311734
rect 274404 276054 275004 311498
rect 274404 275818 274586 276054
rect 274822 275818 275004 276054
rect 274404 275734 275004 275818
rect 274404 275498 274586 275734
rect 274822 275498 275004 275734
rect 274404 240054 275004 275498
rect 274404 239818 274586 240054
rect 274822 239818 275004 240054
rect 274404 239734 275004 239818
rect 274404 239498 274586 239734
rect 274822 239498 275004 239734
rect 274404 204054 275004 239498
rect 274404 203818 274586 204054
rect 274822 203818 275004 204054
rect 274404 203734 275004 203818
rect 274404 203498 274586 203734
rect 274822 203498 275004 203734
rect 274404 168054 275004 203498
rect 274404 167818 274586 168054
rect 274822 167818 275004 168054
rect 274404 167734 275004 167818
rect 274404 167498 274586 167734
rect 274822 167498 275004 167734
rect 274404 132054 275004 167498
rect 274404 131818 274586 132054
rect 274822 131818 275004 132054
rect 274404 131734 275004 131818
rect 274404 131498 274586 131734
rect 274822 131498 275004 131734
rect 274404 96054 275004 131498
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 278004 675654 278604 708882
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 278004 531654 278604 567098
rect 278004 531418 278186 531654
rect 278422 531418 278604 531654
rect 278004 531334 278604 531418
rect 278004 531098 278186 531334
rect 278422 531098 278604 531334
rect 278004 495654 278604 531098
rect 278004 495418 278186 495654
rect 278422 495418 278604 495654
rect 278004 495334 278604 495418
rect 278004 495098 278186 495334
rect 278422 495098 278604 495334
rect 278004 459654 278604 495098
rect 278004 459418 278186 459654
rect 278422 459418 278604 459654
rect 278004 459334 278604 459418
rect 278004 459098 278186 459334
rect 278422 459098 278604 459334
rect 278004 423654 278604 459098
rect 278004 423418 278186 423654
rect 278422 423418 278604 423654
rect 278004 423334 278604 423418
rect 278004 423098 278186 423334
rect 278422 423098 278604 423334
rect 278004 387654 278604 423098
rect 278004 387418 278186 387654
rect 278422 387418 278604 387654
rect 278004 387334 278604 387418
rect 278004 387098 278186 387334
rect 278422 387098 278604 387334
rect 278004 351654 278604 387098
rect 278004 351418 278186 351654
rect 278422 351418 278604 351654
rect 278004 351334 278604 351418
rect 278004 351098 278186 351334
rect 278422 351098 278604 351334
rect 278004 315654 278604 351098
rect 278004 315418 278186 315654
rect 278422 315418 278604 315654
rect 278004 315334 278604 315418
rect 278004 315098 278186 315334
rect 278422 315098 278604 315334
rect 278004 279654 278604 315098
rect 278004 279418 278186 279654
rect 278422 279418 278604 279654
rect 278004 279334 278604 279418
rect 278004 279098 278186 279334
rect 278422 279098 278604 279334
rect 278004 243654 278604 279098
rect 278004 243418 278186 243654
rect 278422 243418 278604 243654
rect 278004 243334 278604 243418
rect 278004 243098 278186 243334
rect 278422 243098 278604 243334
rect 278004 207654 278604 243098
rect 278004 207418 278186 207654
rect 278422 207418 278604 207654
rect 278004 207334 278604 207418
rect 278004 207098 278186 207334
rect 278422 207098 278604 207334
rect 278004 171654 278604 207098
rect 278004 171418 278186 171654
rect 278422 171418 278604 171654
rect 278004 171334 278604 171418
rect 278004 171098 278186 171334
rect 278422 171098 278604 171334
rect 278004 135654 278604 171098
rect 278004 135418 278186 135654
rect 278422 135418 278604 135654
rect 278004 135334 278604 135418
rect 278004 135098 278186 135334
rect 278422 135098 278604 135334
rect 278004 99654 278604 135098
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 277163 63612 277229 63613
rect 277163 63548 277164 63612
rect 277228 63548 277229 63612
rect 277163 63547 277229 63548
rect 277166 63205 277226 63547
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 277163 63204 277229 63205
rect 277163 63140 277164 63204
rect 277228 63140 277229 63204
rect 277163 63139 277229 63140
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 277163 40492 277229 40493
rect 277163 40428 277164 40492
rect 277228 40428 277229 40492
rect 277163 40427 277229 40428
rect 277166 40085 277226 40427
rect 277163 40084 277229 40085
rect 277163 40020 277164 40084
rect 277228 40020 277229 40084
rect 277163 40019 277229 40020
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3106 275004 23498
rect 274404 -3342 274586 -3106
rect 274822 -3342 275004 -3106
rect 274404 -3426 275004 -3342
rect 274404 -3662 274586 -3426
rect 274822 -3662 275004 -3426
rect 274404 -3684 275004 -3662
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -4946 278604 27098
rect 278004 -5182 278186 -4946
rect 278422 -5182 278604 -4946
rect 278004 -5266 278604 -5182
rect 278004 -5502 278186 -5266
rect 278422 -5502 278604 -5266
rect 278004 -5524 278604 -5502
rect 281604 679254 282204 710722
rect 299604 710358 300204 711300
rect 299604 710122 299786 710358
rect 300022 710122 300204 710358
rect 299604 710038 300204 710122
rect 299604 709802 299786 710038
rect 300022 709802 300204 710038
rect 296004 708518 296604 709460
rect 296004 708282 296186 708518
rect 296422 708282 296604 708518
rect 296004 708198 296604 708282
rect 296004 707962 296186 708198
rect 296422 707962 296604 708198
rect 292404 706678 293004 707620
rect 292404 706442 292586 706678
rect 292822 706442 293004 706678
rect 292404 706358 293004 706442
rect 292404 706122 292586 706358
rect 292822 706122 293004 706358
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 281604 535254 282204 570698
rect 281604 535018 281786 535254
rect 282022 535018 282204 535254
rect 281604 534934 282204 535018
rect 281604 534698 281786 534934
rect 282022 534698 282204 534934
rect 281604 499254 282204 534698
rect 281604 499018 281786 499254
rect 282022 499018 282204 499254
rect 281604 498934 282204 499018
rect 281604 498698 281786 498934
rect 282022 498698 282204 498934
rect 281604 463254 282204 498698
rect 281604 463018 281786 463254
rect 282022 463018 282204 463254
rect 281604 462934 282204 463018
rect 281604 462698 281786 462934
rect 282022 462698 282204 462934
rect 281604 427254 282204 462698
rect 281604 427018 281786 427254
rect 282022 427018 282204 427254
rect 281604 426934 282204 427018
rect 281604 426698 281786 426934
rect 282022 426698 282204 426934
rect 281604 391254 282204 426698
rect 281604 391018 281786 391254
rect 282022 391018 282204 391254
rect 281604 390934 282204 391018
rect 281604 390698 281786 390934
rect 282022 390698 282204 390934
rect 281604 355254 282204 390698
rect 281604 355018 281786 355254
rect 282022 355018 282204 355254
rect 281604 354934 282204 355018
rect 281604 354698 281786 354934
rect 282022 354698 282204 354934
rect 281604 319254 282204 354698
rect 281604 319018 281786 319254
rect 282022 319018 282204 319254
rect 281604 318934 282204 319018
rect 281604 318698 281786 318934
rect 282022 318698 282204 318934
rect 281604 283254 282204 318698
rect 281604 283018 281786 283254
rect 282022 283018 282204 283254
rect 281604 282934 282204 283018
rect 281604 282698 281786 282934
rect 282022 282698 282204 282934
rect 281604 247254 282204 282698
rect 281604 247018 281786 247254
rect 282022 247018 282204 247254
rect 281604 246934 282204 247018
rect 281604 246698 281786 246934
rect 282022 246698 282204 246934
rect 281604 211254 282204 246698
rect 281604 211018 281786 211254
rect 282022 211018 282204 211254
rect 281604 210934 282204 211018
rect 281604 210698 281786 210934
rect 282022 210698 282204 210934
rect 281604 175254 282204 210698
rect 281604 175018 281786 175254
rect 282022 175018 282204 175254
rect 281604 174934 282204 175018
rect 281604 174698 281786 174934
rect 282022 174698 282204 174934
rect 281604 139254 282204 174698
rect 281604 139018 281786 139254
rect 282022 139018 282204 139254
rect 281604 138934 282204 139018
rect 281604 138698 281786 138934
rect 282022 138698 282204 138934
rect 281604 103254 282204 138698
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6102 263786 -5866
rect 264022 -6102 264204 -5866
rect 263604 -6186 264204 -6102
rect 263604 -6422 263786 -6186
rect 264022 -6422 264204 -6186
rect 263604 -7364 264204 -6422
rect 281604 -6786 282204 30698
rect 288804 704838 289404 705780
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 288804 326454 289404 361898
rect 288804 326218 288986 326454
rect 289222 326218 289404 326454
rect 288804 326134 289404 326218
rect 288804 325898 288986 326134
rect 289222 325898 289404 326134
rect 288804 290454 289404 325898
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 288804 254454 289404 289898
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 288804 218454 289404 253898
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1844 289404 -902
rect 292404 690054 293004 706122
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 474054 293004 509498
rect 292404 473818 292586 474054
rect 292822 473818 293004 474054
rect 292404 473734 293004 473818
rect 292404 473498 292586 473734
rect 292822 473498 293004 473734
rect 292404 438054 293004 473498
rect 292404 437818 292586 438054
rect 292822 437818 293004 438054
rect 292404 437734 293004 437818
rect 292404 437498 292586 437734
rect 292822 437498 293004 437734
rect 292404 402054 293004 437498
rect 292404 401818 292586 402054
rect 292822 401818 293004 402054
rect 292404 401734 293004 401818
rect 292404 401498 292586 401734
rect 292822 401498 293004 401734
rect 292404 366054 293004 401498
rect 292404 365818 292586 366054
rect 292822 365818 293004 366054
rect 292404 365734 293004 365818
rect 292404 365498 292586 365734
rect 292822 365498 293004 365734
rect 292404 330054 293004 365498
rect 292404 329818 292586 330054
rect 292822 329818 293004 330054
rect 292404 329734 293004 329818
rect 292404 329498 292586 329734
rect 292822 329498 293004 329734
rect 292404 294054 293004 329498
rect 292404 293818 292586 294054
rect 292822 293818 293004 294054
rect 292404 293734 293004 293818
rect 292404 293498 292586 293734
rect 292822 293498 293004 293734
rect 292404 258054 293004 293498
rect 292404 257818 292586 258054
rect 292822 257818 293004 258054
rect 292404 257734 293004 257818
rect 292404 257498 292586 257734
rect 292822 257498 293004 257734
rect 292404 222054 293004 257498
rect 292404 221818 292586 222054
rect 292822 221818 293004 222054
rect 292404 221734 293004 221818
rect 292404 221498 292586 221734
rect 292822 221498 293004 221734
rect 292404 186054 293004 221498
rect 292404 185818 292586 186054
rect 292822 185818 293004 186054
rect 292404 185734 293004 185818
rect 292404 185498 292586 185734
rect 292822 185498 293004 185734
rect 292404 150054 293004 185498
rect 292404 149818 292586 150054
rect 292822 149818 293004 150054
rect 292404 149734 293004 149818
rect 292404 149498 292586 149734
rect 292822 149498 293004 149734
rect 292404 114054 293004 149498
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2186 293004 5498
rect 292404 -2422 292586 -2186
rect 292822 -2422 293004 -2186
rect 292404 -2506 293004 -2422
rect 292404 -2742 292586 -2506
rect 292822 -2742 293004 -2506
rect 292404 -3684 293004 -2742
rect 296004 693654 296604 707962
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 549654 296604 585098
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 296004 513654 296604 549098
rect 296004 513418 296186 513654
rect 296422 513418 296604 513654
rect 296004 513334 296604 513418
rect 296004 513098 296186 513334
rect 296422 513098 296604 513334
rect 296004 477654 296604 513098
rect 296004 477418 296186 477654
rect 296422 477418 296604 477654
rect 296004 477334 296604 477418
rect 296004 477098 296186 477334
rect 296422 477098 296604 477334
rect 296004 441654 296604 477098
rect 296004 441418 296186 441654
rect 296422 441418 296604 441654
rect 296004 441334 296604 441418
rect 296004 441098 296186 441334
rect 296422 441098 296604 441334
rect 296004 405654 296604 441098
rect 296004 405418 296186 405654
rect 296422 405418 296604 405654
rect 296004 405334 296604 405418
rect 296004 405098 296186 405334
rect 296422 405098 296604 405334
rect 296004 369654 296604 405098
rect 296004 369418 296186 369654
rect 296422 369418 296604 369654
rect 296004 369334 296604 369418
rect 296004 369098 296186 369334
rect 296422 369098 296604 369334
rect 296004 333654 296604 369098
rect 296004 333418 296186 333654
rect 296422 333418 296604 333654
rect 296004 333334 296604 333418
rect 296004 333098 296186 333334
rect 296422 333098 296604 333334
rect 296004 297654 296604 333098
rect 296004 297418 296186 297654
rect 296422 297418 296604 297654
rect 296004 297334 296604 297418
rect 296004 297098 296186 297334
rect 296422 297098 296604 297334
rect 296004 261654 296604 297098
rect 296004 261418 296186 261654
rect 296422 261418 296604 261654
rect 296004 261334 296604 261418
rect 296004 261098 296186 261334
rect 296422 261098 296604 261334
rect 296004 225654 296604 261098
rect 296004 225418 296186 225654
rect 296422 225418 296604 225654
rect 296004 225334 296604 225418
rect 296004 225098 296186 225334
rect 296422 225098 296604 225334
rect 296004 189654 296604 225098
rect 296004 189418 296186 189654
rect 296422 189418 296604 189654
rect 296004 189334 296604 189418
rect 296004 189098 296186 189334
rect 296422 189098 296604 189334
rect 296004 153654 296604 189098
rect 296004 153418 296186 153654
rect 296422 153418 296604 153654
rect 296004 153334 296604 153418
rect 296004 153098 296186 153334
rect 296422 153098 296604 153334
rect 296004 117654 296604 153098
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4026 296604 9098
rect 296004 -4262 296186 -4026
rect 296422 -4262 296604 -4026
rect 296004 -4346 296604 -4262
rect 296004 -4582 296186 -4346
rect 296422 -4582 296604 -4346
rect 296004 -5524 296604 -4582
rect 299604 697254 300204 709802
rect 317604 711278 318204 711300
rect 317604 711042 317786 711278
rect 318022 711042 318204 711278
rect 317604 710958 318204 711042
rect 317604 710722 317786 710958
rect 318022 710722 318204 710958
rect 314004 709438 314604 709460
rect 314004 709202 314186 709438
rect 314422 709202 314604 709438
rect 314004 709118 314604 709202
rect 314004 708882 314186 709118
rect 314422 708882 314604 709118
rect 310404 707598 311004 707620
rect 310404 707362 310586 707598
rect 310822 707362 311004 707598
rect 310404 707278 311004 707362
rect 310404 707042 310586 707278
rect 310822 707042 311004 707278
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 589254 300204 624698
rect 299604 589018 299786 589254
rect 300022 589018 300204 589254
rect 299604 588934 300204 589018
rect 299604 588698 299786 588934
rect 300022 588698 300204 588934
rect 299604 553254 300204 588698
rect 299604 553018 299786 553254
rect 300022 553018 300204 553254
rect 299604 552934 300204 553018
rect 299604 552698 299786 552934
rect 300022 552698 300204 552934
rect 299604 517254 300204 552698
rect 299604 517018 299786 517254
rect 300022 517018 300204 517254
rect 299604 516934 300204 517018
rect 299604 516698 299786 516934
rect 300022 516698 300204 516934
rect 299604 481254 300204 516698
rect 299604 481018 299786 481254
rect 300022 481018 300204 481254
rect 299604 480934 300204 481018
rect 299604 480698 299786 480934
rect 300022 480698 300204 480934
rect 299604 445254 300204 480698
rect 299604 445018 299786 445254
rect 300022 445018 300204 445254
rect 299604 444934 300204 445018
rect 299604 444698 299786 444934
rect 300022 444698 300204 444934
rect 299604 409254 300204 444698
rect 299604 409018 299786 409254
rect 300022 409018 300204 409254
rect 299604 408934 300204 409018
rect 299604 408698 299786 408934
rect 300022 408698 300204 408934
rect 299604 373254 300204 408698
rect 299604 373018 299786 373254
rect 300022 373018 300204 373254
rect 299604 372934 300204 373018
rect 299604 372698 299786 372934
rect 300022 372698 300204 372934
rect 299604 337254 300204 372698
rect 299604 337018 299786 337254
rect 300022 337018 300204 337254
rect 299604 336934 300204 337018
rect 299604 336698 299786 336934
rect 300022 336698 300204 336934
rect 299604 301254 300204 336698
rect 299604 301018 299786 301254
rect 300022 301018 300204 301254
rect 299604 300934 300204 301018
rect 299604 300698 299786 300934
rect 300022 300698 300204 300934
rect 299604 265254 300204 300698
rect 299604 265018 299786 265254
rect 300022 265018 300204 265254
rect 299604 264934 300204 265018
rect 299604 264698 299786 264934
rect 300022 264698 300204 264934
rect 299604 229254 300204 264698
rect 299604 229018 299786 229254
rect 300022 229018 300204 229254
rect 299604 228934 300204 229018
rect 299604 228698 299786 228934
rect 300022 228698 300204 228934
rect 299604 193254 300204 228698
rect 299604 193018 299786 193254
rect 300022 193018 300204 193254
rect 299604 192934 300204 193018
rect 299604 192698 299786 192934
rect 300022 192698 300204 192934
rect 299604 157254 300204 192698
rect 299604 157018 299786 157254
rect 300022 157018 300204 157254
rect 299604 156934 300204 157018
rect 299604 156698 299786 156934
rect 300022 156698 300204 156934
rect 299604 121254 300204 156698
rect 299604 121018 299786 121254
rect 300022 121018 300204 121254
rect 299604 120934 300204 121018
rect 299604 120698 299786 120934
rect 300022 120698 300204 120934
rect 299604 85254 300204 120698
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 306804 705758 307404 705780
rect 306804 705522 306986 705758
rect 307222 705522 307404 705758
rect 306804 705438 307404 705522
rect 306804 705202 306986 705438
rect 307222 705202 307404 705438
rect 306804 668454 307404 705202
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306804 560454 307404 595898
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 524454 307404 559898
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 380454 307404 415898
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 306804 344454 307404 379898
rect 306804 344218 306986 344454
rect 307222 344218 307404 344454
rect 306804 344134 307404 344218
rect 306804 343898 306986 344134
rect 307222 343898 307404 344134
rect 306804 308454 307404 343898
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 306804 272454 307404 307898
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 306804 236454 307404 271898
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 200454 307404 235898
rect 306804 200218 306986 200454
rect 307222 200218 307404 200454
rect 306804 200134 307404 200218
rect 306804 199898 306986 200134
rect 307222 199898 307404 200134
rect 306804 164454 307404 199898
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 128454 307404 163898
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 306804 92454 307404 127898
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 302003 16284 302069 16285
rect 302003 16220 302004 16284
rect 302068 16220 302069 16284
rect 302003 16219 302069 16220
rect 302006 15605 302066 16219
rect 302003 15604 302069 15605
rect 302003 15540 302004 15604
rect 302068 15540 302069 15604
rect 302003 15539 302069 15540
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7022 281786 -6786
rect 282022 -7022 282204 -6786
rect 281604 -7106 282204 -7022
rect 281604 -7342 281786 -7106
rect 282022 -7342 282204 -7106
rect 281604 -7364 282204 -7342
rect 299604 -5866 300204 12698
rect 306804 -1266 307404 19898
rect 306804 -1502 306986 -1266
rect 307222 -1502 307404 -1266
rect 306804 -1586 307404 -1502
rect 306804 -1822 306986 -1586
rect 307222 -1822 307404 -1586
rect 306804 -1844 307404 -1822
rect 310404 672054 311004 707042
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 600054 311004 635498
rect 310404 599818 310586 600054
rect 310822 599818 311004 600054
rect 310404 599734 311004 599818
rect 310404 599498 310586 599734
rect 310822 599498 311004 599734
rect 310404 564054 311004 599498
rect 310404 563818 310586 564054
rect 310822 563818 311004 564054
rect 310404 563734 311004 563818
rect 310404 563498 310586 563734
rect 310822 563498 311004 563734
rect 310404 528054 311004 563498
rect 310404 527818 310586 528054
rect 310822 527818 311004 528054
rect 310404 527734 311004 527818
rect 310404 527498 310586 527734
rect 310822 527498 311004 527734
rect 310404 492054 311004 527498
rect 310404 491818 310586 492054
rect 310822 491818 311004 492054
rect 310404 491734 311004 491818
rect 310404 491498 310586 491734
rect 310822 491498 311004 491734
rect 310404 456054 311004 491498
rect 310404 455818 310586 456054
rect 310822 455818 311004 456054
rect 310404 455734 311004 455818
rect 310404 455498 310586 455734
rect 310822 455498 311004 455734
rect 310404 420054 311004 455498
rect 310404 419818 310586 420054
rect 310822 419818 311004 420054
rect 310404 419734 311004 419818
rect 310404 419498 310586 419734
rect 310822 419498 311004 419734
rect 310404 384054 311004 419498
rect 310404 383818 310586 384054
rect 310822 383818 311004 384054
rect 310404 383734 311004 383818
rect 310404 383498 310586 383734
rect 310822 383498 311004 383734
rect 310404 348054 311004 383498
rect 310404 347818 310586 348054
rect 310822 347818 311004 348054
rect 310404 347734 311004 347818
rect 310404 347498 310586 347734
rect 310822 347498 311004 347734
rect 310404 312054 311004 347498
rect 310404 311818 310586 312054
rect 310822 311818 311004 312054
rect 310404 311734 311004 311818
rect 310404 311498 310586 311734
rect 310822 311498 311004 311734
rect 310404 276054 311004 311498
rect 310404 275818 310586 276054
rect 310822 275818 311004 276054
rect 310404 275734 311004 275818
rect 310404 275498 310586 275734
rect 310822 275498 311004 275734
rect 310404 240054 311004 275498
rect 310404 239818 310586 240054
rect 310822 239818 311004 240054
rect 310404 239734 311004 239818
rect 310404 239498 310586 239734
rect 310822 239498 311004 239734
rect 310404 204054 311004 239498
rect 310404 203818 310586 204054
rect 310822 203818 311004 204054
rect 310404 203734 311004 203818
rect 310404 203498 310586 203734
rect 310822 203498 311004 203734
rect 310404 168054 311004 203498
rect 310404 167818 310586 168054
rect 310822 167818 311004 168054
rect 310404 167734 311004 167818
rect 310404 167498 310586 167734
rect 310822 167498 311004 167734
rect 310404 132054 311004 167498
rect 310404 131818 310586 132054
rect 310822 131818 311004 132054
rect 310404 131734 311004 131818
rect 310404 131498 310586 131734
rect 310822 131498 311004 131734
rect 310404 96054 311004 131498
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3106 311004 23498
rect 314004 675654 314604 708882
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 639654 314604 675098
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 314004 639334 314604 639418
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 314004 603654 314604 639098
rect 314004 603418 314186 603654
rect 314422 603418 314604 603654
rect 314004 603334 314604 603418
rect 314004 603098 314186 603334
rect 314422 603098 314604 603334
rect 314004 567654 314604 603098
rect 314004 567418 314186 567654
rect 314422 567418 314604 567654
rect 314004 567334 314604 567418
rect 314004 567098 314186 567334
rect 314422 567098 314604 567334
rect 314004 531654 314604 567098
rect 314004 531418 314186 531654
rect 314422 531418 314604 531654
rect 314004 531334 314604 531418
rect 314004 531098 314186 531334
rect 314422 531098 314604 531334
rect 314004 495654 314604 531098
rect 314004 495418 314186 495654
rect 314422 495418 314604 495654
rect 314004 495334 314604 495418
rect 314004 495098 314186 495334
rect 314422 495098 314604 495334
rect 314004 459654 314604 495098
rect 314004 459418 314186 459654
rect 314422 459418 314604 459654
rect 314004 459334 314604 459418
rect 314004 459098 314186 459334
rect 314422 459098 314604 459334
rect 314004 423654 314604 459098
rect 314004 423418 314186 423654
rect 314422 423418 314604 423654
rect 314004 423334 314604 423418
rect 314004 423098 314186 423334
rect 314422 423098 314604 423334
rect 314004 387654 314604 423098
rect 314004 387418 314186 387654
rect 314422 387418 314604 387654
rect 314004 387334 314604 387418
rect 314004 387098 314186 387334
rect 314422 387098 314604 387334
rect 314004 351654 314604 387098
rect 314004 351418 314186 351654
rect 314422 351418 314604 351654
rect 314004 351334 314604 351418
rect 314004 351098 314186 351334
rect 314422 351098 314604 351334
rect 314004 315654 314604 351098
rect 314004 315418 314186 315654
rect 314422 315418 314604 315654
rect 314004 315334 314604 315418
rect 314004 315098 314186 315334
rect 314422 315098 314604 315334
rect 314004 279654 314604 315098
rect 314004 279418 314186 279654
rect 314422 279418 314604 279654
rect 314004 279334 314604 279418
rect 314004 279098 314186 279334
rect 314422 279098 314604 279334
rect 314004 243654 314604 279098
rect 314004 243418 314186 243654
rect 314422 243418 314604 243654
rect 314004 243334 314604 243418
rect 314004 243098 314186 243334
rect 314422 243098 314604 243334
rect 314004 207654 314604 243098
rect 314004 207418 314186 207654
rect 314422 207418 314604 207654
rect 314004 207334 314604 207418
rect 314004 207098 314186 207334
rect 314422 207098 314604 207334
rect 314004 171654 314604 207098
rect 314004 171418 314186 171654
rect 314422 171418 314604 171654
rect 314004 171334 314604 171418
rect 314004 171098 314186 171334
rect 314422 171098 314604 171334
rect 314004 135654 314604 171098
rect 314004 135418 314186 135654
rect 314422 135418 314604 135654
rect 314004 135334 314604 135418
rect 314004 135098 314186 135334
rect 314422 135098 314604 135334
rect 314004 99654 314604 135098
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 317604 679254 318204 710722
rect 335604 710358 336204 711300
rect 335604 710122 335786 710358
rect 336022 710122 336204 710358
rect 335604 710038 336204 710122
rect 335604 709802 335786 710038
rect 336022 709802 336204 710038
rect 332004 708518 332604 709460
rect 332004 708282 332186 708518
rect 332422 708282 332604 708518
rect 332004 708198 332604 708282
rect 332004 707962 332186 708198
rect 332422 707962 332604 708198
rect 328404 706678 329004 707620
rect 328404 706442 328586 706678
rect 328822 706442 329004 706678
rect 328404 706358 329004 706442
rect 328404 706122 328586 706358
rect 328822 706122 329004 706358
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 317604 607254 318204 642698
rect 317604 607018 317786 607254
rect 318022 607018 318204 607254
rect 317604 606934 318204 607018
rect 317604 606698 317786 606934
rect 318022 606698 318204 606934
rect 317604 571254 318204 606698
rect 317604 571018 317786 571254
rect 318022 571018 318204 571254
rect 317604 570934 318204 571018
rect 317604 570698 317786 570934
rect 318022 570698 318204 570934
rect 317604 535254 318204 570698
rect 317604 535018 317786 535254
rect 318022 535018 318204 535254
rect 317604 534934 318204 535018
rect 317604 534698 317786 534934
rect 318022 534698 318204 534934
rect 317604 499254 318204 534698
rect 317604 499018 317786 499254
rect 318022 499018 318204 499254
rect 317604 498934 318204 499018
rect 317604 498698 317786 498934
rect 318022 498698 318204 498934
rect 317604 463254 318204 498698
rect 317604 463018 317786 463254
rect 318022 463018 318204 463254
rect 317604 462934 318204 463018
rect 317604 462698 317786 462934
rect 318022 462698 318204 462934
rect 317604 427254 318204 462698
rect 324804 704838 325404 705780
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 578454 325404 613898
rect 324804 578218 324986 578454
rect 325222 578218 325404 578454
rect 324804 578134 325404 578218
rect 324804 577898 324986 578134
rect 325222 577898 325404 578134
rect 324804 542454 325404 577898
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 324804 506454 325404 541898
rect 324804 506218 324986 506454
rect 325222 506218 325404 506454
rect 324804 506134 325404 506218
rect 324804 505898 324986 506134
rect 325222 505898 325404 506134
rect 324804 470454 325404 505898
rect 324804 470218 324986 470454
rect 325222 470218 325404 470454
rect 324804 470134 325404 470218
rect 324804 469898 324986 470134
rect 325222 469898 325404 470134
rect 324635 459372 324701 459373
rect 324635 459308 324636 459372
rect 324700 459308 324701 459372
rect 324635 459307 324701 459308
rect 324638 457741 324698 459307
rect 324635 457740 324701 457741
rect 324635 457676 324636 457740
rect 324700 457676 324701 457740
rect 324635 457675 324701 457676
rect 317604 427018 317786 427254
rect 318022 427018 318204 427254
rect 317604 426934 318204 427018
rect 317604 426698 317786 426934
rect 318022 426698 318204 426934
rect 317604 391254 318204 426698
rect 317604 391018 317786 391254
rect 318022 391018 318204 391254
rect 317604 390934 318204 391018
rect 317604 390698 317786 390934
rect 318022 390698 318204 390934
rect 317604 355254 318204 390698
rect 317604 355018 317786 355254
rect 318022 355018 318204 355254
rect 317604 354934 318204 355018
rect 317604 354698 317786 354934
rect 318022 354698 318204 354934
rect 317604 319254 318204 354698
rect 317604 319018 317786 319254
rect 318022 319018 318204 319254
rect 317604 318934 318204 319018
rect 317604 318698 317786 318934
rect 318022 318698 318204 318934
rect 317604 283254 318204 318698
rect 317604 283018 317786 283254
rect 318022 283018 318204 283254
rect 317604 282934 318204 283018
rect 317604 282698 317786 282934
rect 318022 282698 318204 282934
rect 317604 247254 318204 282698
rect 317604 247018 317786 247254
rect 318022 247018 318204 247254
rect 317604 246934 318204 247018
rect 317604 246698 317786 246934
rect 318022 246698 318204 246934
rect 317604 211254 318204 246698
rect 317604 211018 317786 211254
rect 318022 211018 318204 211254
rect 317604 210934 318204 211018
rect 317604 210698 317786 210934
rect 318022 210698 318204 210934
rect 317604 175254 318204 210698
rect 317604 175018 317786 175254
rect 318022 175018 318204 175254
rect 317604 174934 318204 175018
rect 317604 174698 317786 174934
rect 318022 174698 318204 174934
rect 317604 139254 318204 174698
rect 317604 139018 317786 139254
rect 318022 139018 318204 139254
rect 317604 138934 318204 139018
rect 317604 138698 317786 138934
rect 318022 138698 318204 138934
rect 317604 103254 318204 138698
rect 317604 103018 317786 103254
rect 318022 103018 318204 103254
rect 317604 102934 318204 103018
rect 317604 102698 317786 102934
rect 318022 102698 318204 102934
rect 317604 67254 318204 102698
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 315987 63748 316053 63749
rect 315987 63684 315988 63748
rect 316052 63684 316053 63748
rect 315987 63683 316053 63684
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 315990 63341 316050 63683
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 315987 63340 316053 63341
rect 315987 63276 315988 63340
rect 316052 63276 316053 63340
rect 315987 63275 316053 63276
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 313043 16284 313109 16285
rect 313043 16220 313044 16284
rect 313108 16220 313109 16284
rect 313043 16219 313109 16220
rect 313046 15605 313106 16219
rect 313043 15604 313109 15605
rect 313043 15540 313044 15604
rect 313108 15540 313109 15604
rect 313043 15539 313109 15540
rect 310404 -3342 310586 -3106
rect 310822 -3342 311004 -3106
rect 310404 -3426 311004 -3342
rect 310404 -3662 310586 -3426
rect 310822 -3662 311004 -3426
rect 310404 -3684 311004 -3662
rect 314004 -4946 314604 27098
rect 314004 -5182 314186 -4946
rect 314422 -5182 314604 -4946
rect 314004 -5266 314604 -5182
rect 314004 -5502 314186 -5266
rect 314422 -5502 314604 -5266
rect 314004 -5524 314604 -5502
rect 317604 31254 318204 66698
rect 324804 434454 325404 469898
rect 324804 434218 324986 434454
rect 325222 434218 325404 434454
rect 324804 434134 325404 434218
rect 324804 433898 324986 434134
rect 325222 433898 325404 434134
rect 324804 398454 325404 433898
rect 324804 398218 324986 398454
rect 325222 398218 325404 398454
rect 324804 398134 325404 398218
rect 324804 397898 324986 398134
rect 325222 397898 325404 398134
rect 324804 362454 325404 397898
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 324804 290454 325404 325898
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 324804 254454 325404 289898
rect 324804 254218 324986 254454
rect 325222 254218 325404 254454
rect 324804 254134 325404 254218
rect 324804 253898 324986 254134
rect 325222 253898 325404 254134
rect 324804 218454 325404 253898
rect 324804 218218 324986 218454
rect 325222 218218 325404 218454
rect 324804 218134 325404 218218
rect 324804 217898 324986 218134
rect 325222 217898 325404 218134
rect 324804 182454 325404 217898
rect 324804 182218 324986 182454
rect 325222 182218 325404 182454
rect 324804 182134 325404 182218
rect 324804 181898 324986 182134
rect 325222 181898 325404 182134
rect 324804 146454 325404 181898
rect 324804 146218 324986 146454
rect 325222 146218 325404 146454
rect 324804 146134 325404 146218
rect 324804 145898 324986 146134
rect 325222 145898 325404 146134
rect 324804 110454 325404 145898
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 324804 74454 325404 109898
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324267 64020 324333 64021
rect 324267 63956 324268 64020
rect 324332 63956 324333 64020
rect 324267 63955 324333 63956
rect 324270 63749 324330 63955
rect 324267 63748 324333 63749
rect 324267 63684 324268 63748
rect 324332 63684 324333 63748
rect 324267 63683 324333 63684
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6102 299786 -5866
rect 300022 -6102 300204 -5866
rect 299604 -6186 300204 -6102
rect 299604 -6422 299786 -6186
rect 300022 -6422 300204 -6186
rect 299604 -7364 300204 -6422
rect 317604 -6786 318204 30698
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324451 18052 324517 18053
rect 324451 17988 324452 18052
rect 324516 17988 324517 18052
rect 324451 17987 324517 17988
rect 324267 16556 324333 16557
rect 324267 16492 324268 16556
rect 324332 16492 324333 16556
rect 324267 16491 324333 16492
rect 324270 16010 324330 16491
rect 324454 16010 324514 17987
rect 324270 15950 324514 16010
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1844 325404 -902
rect 328404 690054 329004 706122
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 582054 329004 617498
rect 328404 581818 328586 582054
rect 328822 581818 329004 582054
rect 328404 581734 329004 581818
rect 328404 581498 328586 581734
rect 328822 581498 329004 581734
rect 328404 546054 329004 581498
rect 328404 545818 328586 546054
rect 328822 545818 329004 546054
rect 328404 545734 329004 545818
rect 328404 545498 328586 545734
rect 328822 545498 329004 545734
rect 328404 510054 329004 545498
rect 328404 509818 328586 510054
rect 328822 509818 329004 510054
rect 328404 509734 329004 509818
rect 328404 509498 328586 509734
rect 328822 509498 329004 509734
rect 328404 474054 329004 509498
rect 328404 473818 328586 474054
rect 328822 473818 329004 474054
rect 328404 473734 329004 473818
rect 328404 473498 328586 473734
rect 328822 473498 329004 473734
rect 328404 438054 329004 473498
rect 328404 437818 328586 438054
rect 328822 437818 329004 438054
rect 328404 437734 329004 437818
rect 328404 437498 328586 437734
rect 328822 437498 329004 437734
rect 328404 402054 329004 437498
rect 328404 401818 328586 402054
rect 328822 401818 329004 402054
rect 328404 401734 329004 401818
rect 328404 401498 328586 401734
rect 328822 401498 329004 401734
rect 328404 366054 329004 401498
rect 328404 365818 328586 366054
rect 328822 365818 329004 366054
rect 328404 365734 329004 365818
rect 328404 365498 328586 365734
rect 328822 365498 329004 365734
rect 328404 330054 329004 365498
rect 328404 329818 328586 330054
rect 328822 329818 329004 330054
rect 328404 329734 329004 329818
rect 328404 329498 328586 329734
rect 328822 329498 329004 329734
rect 328404 294054 329004 329498
rect 328404 293818 328586 294054
rect 328822 293818 329004 294054
rect 328404 293734 329004 293818
rect 328404 293498 328586 293734
rect 328822 293498 329004 293734
rect 328404 258054 329004 293498
rect 328404 257818 328586 258054
rect 328822 257818 329004 258054
rect 328404 257734 329004 257818
rect 328404 257498 328586 257734
rect 328822 257498 329004 257734
rect 328404 222054 329004 257498
rect 328404 221818 328586 222054
rect 328822 221818 329004 222054
rect 328404 221734 329004 221818
rect 328404 221498 328586 221734
rect 328822 221498 329004 221734
rect 328404 186054 329004 221498
rect 328404 185818 328586 186054
rect 328822 185818 329004 186054
rect 328404 185734 329004 185818
rect 328404 185498 328586 185734
rect 328822 185498 329004 185734
rect 328404 150054 329004 185498
rect 328404 149818 328586 150054
rect 328822 149818 329004 150054
rect 328404 149734 329004 149818
rect 328404 149498 328586 149734
rect 328822 149498 329004 149734
rect 328404 114054 329004 149498
rect 328404 113818 328586 114054
rect 328822 113818 329004 114054
rect 328404 113734 329004 113818
rect 328404 113498 328586 113734
rect 328822 113498 329004 113734
rect 328404 78054 329004 113498
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2186 329004 5498
rect 328404 -2422 328586 -2186
rect 328822 -2422 329004 -2186
rect 328404 -2506 329004 -2422
rect 328404 -2742 328586 -2506
rect 328822 -2742 329004 -2506
rect 328404 -3684 329004 -2742
rect 332004 693654 332604 707962
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 585654 332604 621098
rect 332004 585418 332186 585654
rect 332422 585418 332604 585654
rect 332004 585334 332604 585418
rect 332004 585098 332186 585334
rect 332422 585098 332604 585334
rect 332004 549654 332604 585098
rect 332004 549418 332186 549654
rect 332422 549418 332604 549654
rect 332004 549334 332604 549418
rect 332004 549098 332186 549334
rect 332422 549098 332604 549334
rect 332004 513654 332604 549098
rect 332004 513418 332186 513654
rect 332422 513418 332604 513654
rect 332004 513334 332604 513418
rect 332004 513098 332186 513334
rect 332422 513098 332604 513334
rect 332004 477654 332604 513098
rect 332004 477418 332186 477654
rect 332422 477418 332604 477654
rect 332004 477334 332604 477418
rect 332004 477098 332186 477334
rect 332422 477098 332604 477334
rect 332004 441654 332604 477098
rect 332004 441418 332186 441654
rect 332422 441418 332604 441654
rect 332004 441334 332604 441418
rect 332004 441098 332186 441334
rect 332422 441098 332604 441334
rect 332004 405654 332604 441098
rect 332004 405418 332186 405654
rect 332422 405418 332604 405654
rect 332004 405334 332604 405418
rect 332004 405098 332186 405334
rect 332422 405098 332604 405334
rect 332004 369654 332604 405098
rect 332004 369418 332186 369654
rect 332422 369418 332604 369654
rect 332004 369334 332604 369418
rect 332004 369098 332186 369334
rect 332422 369098 332604 369334
rect 332004 333654 332604 369098
rect 332004 333418 332186 333654
rect 332422 333418 332604 333654
rect 332004 333334 332604 333418
rect 332004 333098 332186 333334
rect 332422 333098 332604 333334
rect 332004 297654 332604 333098
rect 332004 297418 332186 297654
rect 332422 297418 332604 297654
rect 332004 297334 332604 297418
rect 332004 297098 332186 297334
rect 332422 297098 332604 297334
rect 332004 261654 332604 297098
rect 332004 261418 332186 261654
rect 332422 261418 332604 261654
rect 332004 261334 332604 261418
rect 332004 261098 332186 261334
rect 332422 261098 332604 261334
rect 332004 225654 332604 261098
rect 332004 225418 332186 225654
rect 332422 225418 332604 225654
rect 332004 225334 332604 225418
rect 332004 225098 332186 225334
rect 332422 225098 332604 225334
rect 332004 189654 332604 225098
rect 332004 189418 332186 189654
rect 332422 189418 332604 189654
rect 332004 189334 332604 189418
rect 332004 189098 332186 189334
rect 332422 189098 332604 189334
rect 332004 153654 332604 189098
rect 332004 153418 332186 153654
rect 332422 153418 332604 153654
rect 332004 153334 332604 153418
rect 332004 153098 332186 153334
rect 332422 153098 332604 153334
rect 332004 117654 332604 153098
rect 332004 117418 332186 117654
rect 332422 117418 332604 117654
rect 332004 117334 332604 117418
rect 332004 117098 332186 117334
rect 332422 117098 332604 117334
rect 332004 81654 332604 117098
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4026 332604 9098
rect 332004 -4262 332186 -4026
rect 332422 -4262 332604 -4026
rect 332004 -4346 332604 -4262
rect 332004 -4582 332186 -4346
rect 332422 -4582 332604 -4346
rect 332004 -5524 332604 -4582
rect 335604 697254 336204 709802
rect 353604 711278 354204 711300
rect 353604 711042 353786 711278
rect 354022 711042 354204 711278
rect 353604 710958 354204 711042
rect 353604 710722 353786 710958
rect 354022 710722 354204 710958
rect 350004 709438 350604 709460
rect 350004 709202 350186 709438
rect 350422 709202 350604 709438
rect 350004 709118 350604 709202
rect 350004 708882 350186 709118
rect 350422 708882 350604 709118
rect 346404 707598 347004 707620
rect 346404 707362 346586 707598
rect 346822 707362 347004 707598
rect 346404 707278 347004 707362
rect 346404 707042 346586 707278
rect 346822 707042 347004 707278
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 625254 336204 660698
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 589254 336204 624698
rect 335604 589018 335786 589254
rect 336022 589018 336204 589254
rect 335604 588934 336204 589018
rect 335604 588698 335786 588934
rect 336022 588698 336204 588934
rect 335604 553254 336204 588698
rect 335604 553018 335786 553254
rect 336022 553018 336204 553254
rect 335604 552934 336204 553018
rect 335604 552698 335786 552934
rect 336022 552698 336204 552934
rect 335604 517254 336204 552698
rect 335604 517018 335786 517254
rect 336022 517018 336204 517254
rect 335604 516934 336204 517018
rect 335604 516698 335786 516934
rect 336022 516698 336204 516934
rect 335604 481254 336204 516698
rect 335604 481018 335786 481254
rect 336022 481018 336204 481254
rect 335604 480934 336204 481018
rect 335604 480698 335786 480934
rect 336022 480698 336204 480934
rect 335604 445254 336204 480698
rect 342804 705758 343404 705780
rect 342804 705522 342986 705758
rect 343222 705522 343404 705758
rect 342804 705438 343404 705522
rect 342804 705202 342986 705438
rect 343222 705202 343404 705438
rect 342804 668454 343404 705202
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 560454 343404 595898
rect 342804 560218 342986 560454
rect 343222 560218 343404 560454
rect 342804 560134 343404 560218
rect 342804 559898 342986 560134
rect 343222 559898 343404 560134
rect 342804 524454 343404 559898
rect 342804 524218 342986 524454
rect 343222 524218 343404 524454
rect 342804 524134 343404 524218
rect 342804 523898 342986 524134
rect 343222 523898 343404 524134
rect 342804 488454 343404 523898
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342483 459780 342549 459781
rect 342483 459716 342484 459780
rect 342548 459716 342549 459780
rect 342483 459715 342549 459716
rect 335604 445018 335786 445254
rect 336022 445018 336204 445254
rect 335604 444934 336204 445018
rect 335604 444698 335786 444934
rect 336022 444698 336204 444934
rect 335604 409254 336204 444698
rect 335604 409018 335786 409254
rect 336022 409018 336204 409254
rect 335604 408934 336204 409018
rect 335604 408698 335786 408934
rect 336022 408698 336204 408934
rect 335604 373254 336204 408698
rect 335604 373018 335786 373254
rect 336022 373018 336204 373254
rect 335604 372934 336204 373018
rect 335604 372698 335786 372934
rect 336022 372698 336204 372934
rect 335604 337254 336204 372698
rect 335604 337018 335786 337254
rect 336022 337018 336204 337254
rect 335604 336934 336204 337018
rect 335604 336698 335786 336934
rect 336022 336698 336204 336934
rect 335604 301254 336204 336698
rect 335604 301018 335786 301254
rect 336022 301018 336204 301254
rect 335604 300934 336204 301018
rect 335604 300698 335786 300934
rect 336022 300698 336204 300934
rect 335604 265254 336204 300698
rect 335604 265018 335786 265254
rect 336022 265018 336204 265254
rect 335604 264934 336204 265018
rect 335604 264698 335786 264934
rect 336022 264698 336204 264934
rect 335604 229254 336204 264698
rect 335604 229018 335786 229254
rect 336022 229018 336204 229254
rect 335604 228934 336204 229018
rect 335604 228698 335786 228934
rect 336022 228698 336204 228934
rect 335604 193254 336204 228698
rect 342486 216885 342546 459715
rect 342667 459644 342733 459645
rect 342667 459580 342668 459644
rect 342732 459580 342733 459644
rect 342667 459579 342733 459580
rect 342483 216884 342549 216885
rect 342483 216820 342484 216884
rect 342548 216820 342549 216884
rect 342483 216819 342549 216820
rect 335604 193018 335786 193254
rect 336022 193018 336204 193254
rect 335604 192934 336204 193018
rect 335604 192698 335786 192934
rect 336022 192698 336204 192934
rect 335604 157254 336204 192698
rect 342670 169965 342730 459579
rect 342804 452454 343404 487898
rect 346404 672054 347004 707042
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 600054 347004 635498
rect 346404 599818 346586 600054
rect 346822 599818 347004 600054
rect 346404 599734 347004 599818
rect 346404 599498 346586 599734
rect 346822 599498 347004 599734
rect 346404 564054 347004 599498
rect 346404 563818 346586 564054
rect 346822 563818 347004 564054
rect 346404 563734 347004 563818
rect 346404 563498 346586 563734
rect 346822 563498 347004 563734
rect 346404 528054 347004 563498
rect 346404 527818 346586 528054
rect 346822 527818 347004 528054
rect 346404 527734 347004 527818
rect 346404 527498 346586 527734
rect 346822 527498 347004 527734
rect 346404 492054 347004 527498
rect 346404 491818 346586 492054
rect 346822 491818 347004 492054
rect 346404 491734 347004 491818
rect 346404 491498 346586 491734
rect 346822 491498 347004 491734
rect 344323 460052 344389 460053
rect 344323 459988 344324 460052
rect 344388 459988 344389 460052
rect 344323 459987 344389 459988
rect 344139 459916 344205 459917
rect 344139 459852 344140 459916
rect 344204 459852 344205 459916
rect 344139 459851 344205 459852
rect 343587 459644 343653 459645
rect 343587 459580 343588 459644
rect 343652 459580 343653 459644
rect 343587 459579 343653 459580
rect 342804 452218 342986 452454
rect 343222 452218 343404 452454
rect 342804 452134 343404 452218
rect 342804 451898 342986 452134
rect 343222 451898 343404 452134
rect 342804 416454 343404 451898
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 380454 343404 415898
rect 342804 380218 342986 380454
rect 343222 380218 343404 380454
rect 342804 380134 343404 380218
rect 342804 379898 342986 380134
rect 343222 379898 343404 380134
rect 342804 344454 343404 379898
rect 342804 344218 342986 344454
rect 343222 344218 343404 344454
rect 342804 344134 343404 344218
rect 342804 343898 342986 344134
rect 343222 343898 343404 344134
rect 342804 308454 343404 343898
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 342804 272454 343404 307898
rect 342804 272218 342986 272454
rect 343222 272218 343404 272454
rect 342804 272134 343404 272218
rect 342804 271898 342986 272134
rect 343222 271898 343404 272134
rect 342804 236454 343404 271898
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 342804 200454 343404 235898
rect 342804 200218 342986 200454
rect 343222 200218 343404 200454
rect 342804 200134 343404 200218
rect 342804 199898 342986 200134
rect 343222 199898 343404 200134
rect 342667 169964 342733 169965
rect 342667 169900 342668 169964
rect 342732 169900 342733 169964
rect 342667 169899 342733 169900
rect 335604 157018 335786 157254
rect 336022 157018 336204 157254
rect 335604 156934 336204 157018
rect 335604 156698 335786 156934
rect 336022 156698 336204 156934
rect 335604 121254 336204 156698
rect 335604 121018 335786 121254
rect 336022 121018 336204 121254
rect 335604 120934 336204 121018
rect 335604 120698 335786 120934
rect 336022 120698 336204 120934
rect 335604 85254 336204 120698
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 342804 164454 343404 199898
rect 342804 164218 342986 164454
rect 343222 164218 343404 164454
rect 342804 164134 343404 164218
rect 342804 163898 342986 164134
rect 343222 163898 343404 164134
rect 342804 128454 343404 163898
rect 342804 128218 342986 128454
rect 343222 128218 343404 128454
rect 342804 128134 343404 128218
rect 342804 127898 342986 128134
rect 343222 127898 343404 128134
rect 342804 92454 343404 127898
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 343590 80069 343650 459579
rect 344142 263805 344202 459851
rect 344326 310725 344386 459987
rect 345427 459644 345493 459645
rect 345427 459580 345428 459644
rect 345492 459580 345493 459644
rect 345427 459579 345493 459580
rect 345243 459372 345309 459373
rect 345243 459308 345244 459372
rect 345308 459308 345309 459372
rect 345243 459307 345309 459308
rect 344323 310724 344389 310725
rect 344323 310660 344324 310724
rect 344388 310660 344389 310724
rect 344323 310659 344389 310660
rect 344139 263804 344205 263805
rect 344139 263740 344140 263804
rect 344204 263740 344205 263804
rect 344139 263739 344205 263740
rect 343587 80068 343653 80069
rect 343587 80004 343588 80068
rect 343652 80004 343653 80068
rect 343587 80003 343653 80004
rect 345246 64837 345306 459307
rect 345243 64836 345309 64837
rect 345243 64772 345244 64836
rect 345308 64772 345309 64836
rect 345243 64771 345309 64772
rect 343587 64020 343653 64021
rect 343587 63956 343588 64020
rect 343652 63956 343653 64020
rect 343587 63955 343653 63956
rect 343590 63749 343650 63955
rect 343587 63748 343653 63749
rect 343587 63684 343588 63748
rect 343652 63684 343653 63748
rect 343587 63683 343653 63684
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 345430 50965 345490 459579
rect 346404 456054 347004 491498
rect 350004 675654 350604 708882
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 639654 350604 675098
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 603654 350604 639098
rect 350004 603418 350186 603654
rect 350422 603418 350604 603654
rect 350004 603334 350604 603418
rect 350004 603098 350186 603334
rect 350422 603098 350604 603334
rect 350004 567654 350604 603098
rect 350004 567418 350186 567654
rect 350422 567418 350604 567654
rect 350004 567334 350604 567418
rect 350004 567098 350186 567334
rect 350422 567098 350604 567334
rect 350004 531654 350604 567098
rect 350004 531418 350186 531654
rect 350422 531418 350604 531654
rect 350004 531334 350604 531418
rect 350004 531098 350186 531334
rect 350422 531098 350604 531334
rect 350004 495654 350604 531098
rect 350004 495418 350186 495654
rect 350422 495418 350604 495654
rect 350004 495334 350604 495418
rect 350004 495098 350186 495334
rect 350422 495098 350604 495334
rect 348371 463044 348437 463045
rect 348371 462980 348372 463044
rect 348436 462980 348437 463044
rect 348371 462979 348437 462980
rect 347083 459372 347149 459373
rect 347083 459308 347084 459372
rect 347148 459308 347149 459372
rect 347083 459307 347149 459308
rect 346404 455818 346586 456054
rect 346822 455818 347004 456054
rect 346404 455734 347004 455818
rect 346404 455498 346586 455734
rect 346822 455498 347004 455734
rect 346404 420054 347004 455498
rect 346404 419818 346586 420054
rect 346822 419818 347004 420054
rect 346404 419734 347004 419818
rect 346404 419498 346586 419734
rect 346822 419498 347004 419734
rect 346404 384054 347004 419498
rect 346404 383818 346586 384054
rect 346822 383818 347004 384054
rect 346404 383734 347004 383818
rect 346404 383498 346586 383734
rect 346822 383498 347004 383734
rect 346404 348054 347004 383498
rect 346404 347818 346586 348054
rect 346822 347818 347004 348054
rect 346404 347734 347004 347818
rect 346404 347498 346586 347734
rect 346822 347498 347004 347734
rect 346404 312054 347004 347498
rect 346404 311818 346586 312054
rect 346822 311818 347004 312054
rect 346404 311734 347004 311818
rect 346404 311498 346586 311734
rect 346822 311498 347004 311734
rect 346404 276054 347004 311498
rect 346404 275818 346586 276054
rect 346822 275818 347004 276054
rect 346404 275734 347004 275818
rect 346404 275498 346586 275734
rect 346822 275498 347004 275734
rect 346404 240054 347004 275498
rect 346404 239818 346586 240054
rect 346822 239818 347004 240054
rect 346404 239734 347004 239818
rect 346404 239498 346586 239734
rect 346822 239498 347004 239734
rect 346404 204054 347004 239498
rect 346404 203818 346586 204054
rect 346822 203818 347004 204054
rect 346404 203734 347004 203818
rect 346404 203498 346586 203734
rect 346822 203498 347004 203734
rect 346404 168054 347004 203498
rect 346404 167818 346586 168054
rect 346822 167818 347004 168054
rect 346404 167734 347004 167818
rect 346404 167498 346586 167734
rect 346822 167498 347004 167734
rect 346404 132054 347004 167498
rect 346404 131818 346586 132054
rect 346822 131818 347004 132054
rect 346404 131734 347004 131818
rect 346404 131498 346586 131734
rect 346822 131498 347004 131734
rect 346404 96054 347004 131498
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 345427 50964 345493 50965
rect 345427 50900 345428 50964
rect 345492 50900 345493 50964
rect 345427 50899 345493 50900
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 336963 16692 337029 16693
rect 336963 16628 336964 16692
rect 337028 16628 337029 16692
rect 336963 16627 337029 16628
rect 336966 16285 337026 16627
rect 336963 16284 337029 16285
rect 336963 16220 336964 16284
rect 337028 16220 337029 16284
rect 336963 16219 337029 16220
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7022 317786 -6786
rect 318022 -7022 318204 -6786
rect 317604 -7106 318204 -7022
rect 317604 -7342 317786 -7106
rect 318022 -7342 318204 -7106
rect 317604 -7364 318204 -7342
rect 335604 -5866 336204 12698
rect 342804 -1266 343404 19898
rect 342804 -1502 342986 -1266
rect 343222 -1502 343404 -1266
rect 342804 -1586 343404 -1502
rect 342804 -1822 342986 -1586
rect 343222 -1822 343404 -1586
rect 342804 -1844 343404 -1822
rect 346404 24054 347004 59498
rect 347086 35869 347146 459307
rect 348374 345405 348434 462979
rect 348739 462772 348805 462773
rect 348739 462708 348740 462772
rect 348804 462708 348805 462772
rect 348739 462707 348805 462708
rect 348555 462500 348621 462501
rect 348555 462436 348556 462500
rect 348620 462436 348621 462500
rect 348555 462435 348621 462436
rect 348558 368797 348618 462435
rect 348742 392325 348802 462707
rect 348923 462636 348989 462637
rect 348923 462572 348924 462636
rect 348988 462572 348989 462636
rect 348923 462571 348989 462572
rect 348926 415717 348986 462571
rect 350004 459654 350604 495098
rect 350004 459418 350186 459654
rect 350422 459418 350604 459654
rect 350004 459334 350604 459418
rect 350004 459098 350186 459334
rect 350422 459098 350604 459334
rect 350004 423654 350604 459098
rect 350004 423418 350186 423654
rect 350422 423418 350604 423654
rect 350004 423334 350604 423418
rect 350004 423098 350186 423334
rect 350422 423098 350604 423334
rect 348923 415716 348989 415717
rect 348923 415652 348924 415716
rect 348988 415652 348989 415716
rect 348923 415651 348989 415652
rect 348739 392324 348805 392325
rect 348739 392260 348740 392324
rect 348804 392260 348805 392324
rect 348739 392259 348805 392260
rect 350004 387654 350604 423098
rect 350004 387418 350186 387654
rect 350422 387418 350604 387654
rect 350004 387334 350604 387418
rect 350004 387098 350186 387334
rect 350422 387098 350604 387334
rect 348555 368796 348621 368797
rect 348555 368732 348556 368796
rect 348620 368732 348621 368796
rect 348555 368731 348621 368732
rect 350004 351654 350604 387098
rect 350004 351418 350186 351654
rect 350422 351418 350604 351654
rect 350004 351334 350604 351418
rect 350004 351098 350186 351334
rect 350422 351098 350604 351334
rect 348371 345404 348437 345405
rect 348371 345340 348372 345404
rect 348436 345340 348437 345404
rect 348371 345339 348437 345340
rect 350004 315654 350604 351098
rect 350004 315418 350186 315654
rect 350422 315418 350604 315654
rect 350004 315334 350604 315418
rect 350004 315098 350186 315334
rect 350422 315098 350604 315334
rect 350004 279654 350604 315098
rect 350004 279418 350186 279654
rect 350422 279418 350604 279654
rect 350004 279334 350604 279418
rect 350004 279098 350186 279334
rect 350422 279098 350604 279334
rect 350004 243654 350604 279098
rect 350004 243418 350186 243654
rect 350422 243418 350604 243654
rect 350004 243334 350604 243418
rect 350004 243098 350186 243334
rect 350422 243098 350604 243334
rect 350004 207654 350604 243098
rect 350004 207418 350186 207654
rect 350422 207418 350604 207654
rect 350004 207334 350604 207418
rect 350004 207098 350186 207334
rect 350422 207098 350604 207334
rect 350004 171654 350604 207098
rect 350004 171418 350186 171654
rect 350422 171418 350604 171654
rect 350004 171334 350604 171418
rect 350004 171098 350186 171334
rect 350422 171098 350604 171334
rect 350004 135654 350604 171098
rect 350004 135418 350186 135654
rect 350422 135418 350604 135654
rect 350004 135334 350604 135418
rect 350004 135098 350186 135334
rect 350422 135098 350604 135334
rect 350004 99654 350604 135098
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 347083 35868 347149 35869
rect 347083 35804 347084 35868
rect 347148 35804 347149 35868
rect 347083 35803 347149 35804
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3106 347004 23498
rect 346404 -3342 346586 -3106
rect 346822 -3342 347004 -3106
rect 346404 -3426 347004 -3342
rect 346404 -3662 346586 -3426
rect 346822 -3662 347004 -3426
rect 346404 -3684 347004 -3662
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -4946 350604 27098
rect 350004 -5182 350186 -4946
rect 350422 -5182 350604 -4946
rect 350004 -5266 350604 -5182
rect 350004 -5502 350186 -5266
rect 350422 -5502 350604 -5266
rect 350004 -5524 350604 -5502
rect 353604 679254 354204 710722
rect 371604 710358 372204 711300
rect 371604 710122 371786 710358
rect 372022 710122 372204 710358
rect 371604 710038 372204 710122
rect 371604 709802 371786 710038
rect 372022 709802 372204 710038
rect 368004 708518 368604 709460
rect 368004 708282 368186 708518
rect 368422 708282 368604 708518
rect 368004 708198 368604 708282
rect 368004 707962 368186 708198
rect 368422 707962 368604 708198
rect 364404 706678 365004 707620
rect 364404 706442 364586 706678
rect 364822 706442 365004 706678
rect 364404 706358 365004 706442
rect 364404 706122 364586 706358
rect 364822 706122 365004 706358
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 353604 607254 354204 642698
rect 353604 607018 353786 607254
rect 354022 607018 354204 607254
rect 353604 606934 354204 607018
rect 353604 606698 353786 606934
rect 354022 606698 354204 606934
rect 353604 571254 354204 606698
rect 353604 571018 353786 571254
rect 354022 571018 354204 571254
rect 353604 570934 354204 571018
rect 353604 570698 353786 570934
rect 354022 570698 354204 570934
rect 353604 535254 354204 570698
rect 353604 535018 353786 535254
rect 354022 535018 354204 535254
rect 353604 534934 354204 535018
rect 353604 534698 353786 534934
rect 354022 534698 354204 534934
rect 353604 499254 354204 534698
rect 353604 499018 353786 499254
rect 354022 499018 354204 499254
rect 353604 498934 354204 499018
rect 353604 498698 353786 498934
rect 354022 498698 354204 498934
rect 353604 463254 354204 498698
rect 353604 463018 353786 463254
rect 354022 463018 354204 463254
rect 353604 462934 354204 463018
rect 353604 462698 353786 462934
rect 354022 462698 354204 462934
rect 353604 427254 354204 462698
rect 353604 427018 353786 427254
rect 354022 427018 354204 427254
rect 353604 426934 354204 427018
rect 353604 426698 353786 426934
rect 354022 426698 354204 426934
rect 353604 391254 354204 426698
rect 353604 391018 353786 391254
rect 354022 391018 354204 391254
rect 353604 390934 354204 391018
rect 353604 390698 353786 390934
rect 354022 390698 354204 390934
rect 353604 355254 354204 390698
rect 353604 355018 353786 355254
rect 354022 355018 354204 355254
rect 353604 354934 354204 355018
rect 353604 354698 353786 354934
rect 354022 354698 354204 354934
rect 353604 319254 354204 354698
rect 353604 319018 353786 319254
rect 354022 319018 354204 319254
rect 353604 318934 354204 319018
rect 353604 318698 353786 318934
rect 354022 318698 354204 318934
rect 353604 283254 354204 318698
rect 360804 704838 361404 705780
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 578454 361404 613898
rect 360804 578218 360986 578454
rect 361222 578218 361404 578454
rect 360804 578134 361404 578218
rect 360804 577898 360986 578134
rect 361222 577898 361404 578134
rect 360804 542454 361404 577898
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 360804 506454 361404 541898
rect 360804 506218 360986 506454
rect 361222 506218 361404 506454
rect 360804 506134 361404 506218
rect 360804 505898 360986 506134
rect 361222 505898 361404 506134
rect 360804 470454 361404 505898
rect 360804 470218 360986 470454
rect 361222 470218 361404 470454
rect 360804 470134 361404 470218
rect 360804 469898 360986 470134
rect 361222 469898 361404 470134
rect 360804 434454 361404 469898
rect 360804 434218 360986 434454
rect 361222 434218 361404 434454
rect 360804 434134 361404 434218
rect 360804 433898 360986 434134
rect 361222 433898 361404 434134
rect 360804 398454 361404 433898
rect 360804 398218 360986 398454
rect 361222 398218 361404 398454
rect 360804 398134 361404 398218
rect 360804 397898 360986 398134
rect 361222 397898 361404 398134
rect 360804 362454 361404 397898
rect 360804 362218 360986 362454
rect 361222 362218 361404 362454
rect 360804 362134 361404 362218
rect 360804 361898 360986 362134
rect 361222 361898 361404 362134
rect 360804 326454 361404 361898
rect 360804 326218 360986 326454
rect 361222 326218 361404 326454
rect 360804 326134 361404 326218
rect 360804 325898 360986 326134
rect 361222 325898 361404 326134
rect 357387 310588 357453 310589
rect 357387 310524 357388 310588
rect 357452 310524 357453 310588
rect 357387 310523 357453 310524
rect 357390 310317 357450 310523
rect 357387 310316 357453 310317
rect 357387 310252 357388 310316
rect 357452 310252 357453 310316
rect 357387 310251 357453 310252
rect 353604 283018 353786 283254
rect 354022 283018 354204 283254
rect 353604 282934 354204 283018
rect 353604 282698 353786 282934
rect 354022 282698 354204 282934
rect 353604 247254 354204 282698
rect 360804 290454 361404 325898
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 357387 263668 357453 263669
rect 357387 263604 357388 263668
rect 357452 263604 357453 263668
rect 357387 263603 357453 263604
rect 357390 263397 357450 263603
rect 357387 263396 357453 263397
rect 357387 263332 357388 263396
rect 357452 263332 357453 263396
rect 357387 263331 357453 263332
rect 353604 247018 353786 247254
rect 354022 247018 354204 247254
rect 353604 246934 354204 247018
rect 353604 246698 353786 246934
rect 354022 246698 354204 246934
rect 353604 211254 354204 246698
rect 360804 254454 361404 289898
rect 360804 254218 360986 254454
rect 361222 254218 361404 254454
rect 360804 254134 361404 254218
rect 360804 253898 360986 254134
rect 361222 253898 361404 254134
rect 360804 218454 361404 253898
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 357387 216748 357453 216749
rect 357387 216684 357388 216748
rect 357452 216684 357453 216748
rect 357387 216683 357453 216684
rect 357390 216477 357450 216683
rect 357387 216476 357453 216477
rect 357387 216412 357388 216476
rect 357452 216412 357453 216476
rect 357387 216411 357453 216412
rect 353604 211018 353786 211254
rect 354022 211018 354204 211254
rect 353604 210934 354204 211018
rect 353604 210698 353786 210934
rect 354022 210698 354204 210934
rect 353604 175254 354204 210698
rect 353604 175018 353786 175254
rect 354022 175018 354204 175254
rect 353604 174934 354204 175018
rect 353604 174698 353786 174934
rect 354022 174698 354204 174934
rect 353604 139254 354204 174698
rect 360804 182454 361404 217898
rect 360804 182218 360986 182454
rect 361222 182218 361404 182454
rect 360804 182134 361404 182218
rect 360804 181898 360986 182134
rect 361222 181898 361404 182134
rect 357387 169828 357453 169829
rect 357387 169764 357388 169828
rect 357452 169764 357453 169828
rect 357387 169763 357453 169764
rect 357390 169557 357450 169763
rect 357387 169556 357453 169557
rect 357387 169492 357388 169556
rect 357452 169492 357453 169556
rect 357387 169491 357453 169492
rect 353604 139018 353786 139254
rect 354022 139018 354204 139254
rect 353604 138934 354204 139018
rect 353604 138698 353786 138934
rect 354022 138698 354204 138934
rect 353604 103254 354204 138698
rect 353604 103018 353786 103254
rect 354022 103018 354204 103254
rect 353604 102934 354204 103018
rect 353604 102698 353786 102934
rect 354022 102698 354204 102934
rect 353604 67254 354204 102698
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 360804 146454 361404 181898
rect 360804 146218 360986 146454
rect 361222 146218 361404 146454
rect 360804 146134 361404 146218
rect 360804 145898 360986 146134
rect 361222 145898 361404 146134
rect 360804 110454 361404 145898
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 357387 40084 357453 40085
rect 357387 40020 357388 40084
rect 357452 40020 357453 40084
rect 357387 40019 357453 40020
rect 357390 39813 357450 40019
rect 357387 39812 357453 39813
rect 357387 39748 357388 39812
rect 357452 39748 357453 39812
rect 357387 39747 357453 39748
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6102 335786 -5866
rect 336022 -6102 336204 -5866
rect 335604 -6186 336204 -6102
rect 335604 -6422 335786 -6186
rect 336022 -6422 336204 -6186
rect 335604 -7364 336204 -6422
rect 353604 -6786 354204 30698
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1844 361404 -902
rect 364404 690054 365004 706122
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 582054 365004 617498
rect 364404 581818 364586 582054
rect 364822 581818 365004 582054
rect 364404 581734 365004 581818
rect 364404 581498 364586 581734
rect 364822 581498 365004 581734
rect 364404 546054 365004 581498
rect 364404 545818 364586 546054
rect 364822 545818 365004 546054
rect 364404 545734 365004 545818
rect 364404 545498 364586 545734
rect 364822 545498 365004 545734
rect 364404 510054 365004 545498
rect 364404 509818 364586 510054
rect 364822 509818 365004 510054
rect 364404 509734 365004 509818
rect 364404 509498 364586 509734
rect 364822 509498 365004 509734
rect 364404 474054 365004 509498
rect 364404 473818 364586 474054
rect 364822 473818 365004 474054
rect 364404 473734 365004 473818
rect 364404 473498 364586 473734
rect 364822 473498 365004 473734
rect 364404 438054 365004 473498
rect 364404 437818 364586 438054
rect 364822 437818 365004 438054
rect 364404 437734 365004 437818
rect 364404 437498 364586 437734
rect 364822 437498 365004 437734
rect 364404 402054 365004 437498
rect 364404 401818 364586 402054
rect 364822 401818 365004 402054
rect 364404 401734 365004 401818
rect 364404 401498 364586 401734
rect 364822 401498 365004 401734
rect 364404 366054 365004 401498
rect 364404 365818 364586 366054
rect 364822 365818 365004 366054
rect 364404 365734 365004 365818
rect 364404 365498 364586 365734
rect 364822 365498 365004 365734
rect 364404 330054 365004 365498
rect 364404 329818 364586 330054
rect 364822 329818 365004 330054
rect 364404 329734 365004 329818
rect 364404 329498 364586 329734
rect 364822 329498 365004 329734
rect 364404 294054 365004 329498
rect 364404 293818 364586 294054
rect 364822 293818 365004 294054
rect 364404 293734 365004 293818
rect 364404 293498 364586 293734
rect 364822 293498 365004 293734
rect 364404 258054 365004 293498
rect 364404 257818 364586 258054
rect 364822 257818 365004 258054
rect 364404 257734 365004 257818
rect 364404 257498 364586 257734
rect 364822 257498 365004 257734
rect 364404 222054 365004 257498
rect 364404 221818 364586 222054
rect 364822 221818 365004 222054
rect 364404 221734 365004 221818
rect 364404 221498 364586 221734
rect 364822 221498 365004 221734
rect 364404 186054 365004 221498
rect 364404 185818 364586 186054
rect 364822 185818 365004 186054
rect 364404 185734 365004 185818
rect 364404 185498 364586 185734
rect 364822 185498 365004 185734
rect 364404 150054 365004 185498
rect 364404 149818 364586 150054
rect 364822 149818 365004 150054
rect 364404 149734 365004 149818
rect 364404 149498 364586 149734
rect 364822 149498 365004 149734
rect 364404 114054 365004 149498
rect 364404 113818 364586 114054
rect 364822 113818 365004 114054
rect 364404 113734 365004 113818
rect 364404 113498 364586 113734
rect 364822 113498 365004 113734
rect 364404 78054 365004 113498
rect 368004 693654 368604 707962
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 621654 368604 657098
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 585654 368604 621098
rect 368004 585418 368186 585654
rect 368422 585418 368604 585654
rect 368004 585334 368604 585418
rect 368004 585098 368186 585334
rect 368422 585098 368604 585334
rect 368004 549654 368604 585098
rect 368004 549418 368186 549654
rect 368422 549418 368604 549654
rect 368004 549334 368604 549418
rect 368004 549098 368186 549334
rect 368422 549098 368604 549334
rect 368004 513654 368604 549098
rect 368004 513418 368186 513654
rect 368422 513418 368604 513654
rect 368004 513334 368604 513418
rect 368004 513098 368186 513334
rect 368422 513098 368604 513334
rect 368004 477654 368604 513098
rect 368004 477418 368186 477654
rect 368422 477418 368604 477654
rect 368004 477334 368604 477418
rect 368004 477098 368186 477334
rect 368422 477098 368604 477334
rect 368004 441654 368604 477098
rect 368004 441418 368186 441654
rect 368422 441418 368604 441654
rect 368004 441334 368604 441418
rect 368004 441098 368186 441334
rect 368422 441098 368604 441334
rect 368004 405654 368604 441098
rect 368004 405418 368186 405654
rect 368422 405418 368604 405654
rect 368004 405334 368604 405418
rect 368004 405098 368186 405334
rect 368422 405098 368604 405334
rect 368004 369654 368604 405098
rect 368004 369418 368186 369654
rect 368422 369418 368604 369654
rect 368004 369334 368604 369418
rect 368004 369098 368186 369334
rect 368422 369098 368604 369334
rect 368004 333654 368604 369098
rect 368004 333418 368186 333654
rect 368422 333418 368604 333654
rect 368004 333334 368604 333418
rect 368004 333098 368186 333334
rect 368422 333098 368604 333334
rect 368004 297654 368604 333098
rect 368004 297418 368186 297654
rect 368422 297418 368604 297654
rect 368004 297334 368604 297418
rect 368004 297098 368186 297334
rect 368422 297098 368604 297334
rect 368004 261654 368604 297098
rect 368004 261418 368186 261654
rect 368422 261418 368604 261654
rect 368004 261334 368604 261418
rect 368004 261098 368186 261334
rect 368422 261098 368604 261334
rect 368004 225654 368604 261098
rect 368004 225418 368186 225654
rect 368422 225418 368604 225654
rect 368004 225334 368604 225418
rect 368004 225098 368186 225334
rect 368422 225098 368604 225334
rect 368004 189654 368604 225098
rect 368004 189418 368186 189654
rect 368422 189418 368604 189654
rect 368004 189334 368604 189418
rect 368004 189098 368186 189334
rect 368422 189098 368604 189334
rect 368004 153654 368604 189098
rect 368004 153418 368186 153654
rect 368422 153418 368604 153654
rect 368004 153334 368604 153418
rect 368004 153098 368186 153334
rect 368422 153098 368604 153334
rect 368004 117654 368604 153098
rect 368004 117418 368186 117654
rect 368422 117418 368604 117654
rect 368004 117334 368604 117418
rect 368004 117098 368186 117334
rect 368422 117098 368604 117334
rect 365667 87412 365733 87413
rect 365667 87348 365668 87412
rect 365732 87348 365733 87412
rect 365667 87347 365733 87348
rect 365670 87141 365730 87347
rect 365667 87140 365733 87141
rect 365667 87076 365668 87140
rect 365732 87076 365733 87140
rect 365667 87075 365733 87076
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 368004 81654 368604 117098
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 365667 29476 365733 29477
rect 365667 29412 365668 29476
rect 365732 29412 365733 29476
rect 365667 29411 365733 29412
rect 365670 29205 365730 29411
rect 365667 29204 365733 29205
rect 365667 29140 365668 29204
rect 365732 29140 365733 29204
rect 365667 29139 365733 29140
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2186 365004 5498
rect 364404 -2422 364586 -2186
rect 364822 -2422 365004 -2186
rect 364404 -2506 365004 -2422
rect 364404 -2742 364586 -2506
rect 364822 -2742 365004 -2506
rect 364404 -3684 365004 -2742
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4026 368604 9098
rect 368004 -4262 368186 -4026
rect 368422 -4262 368604 -4026
rect 368004 -4346 368604 -4262
rect 368004 -4582 368186 -4346
rect 368422 -4582 368604 -4346
rect 368004 -5524 368604 -4582
rect 371604 697254 372204 709802
rect 389604 711278 390204 711300
rect 389604 711042 389786 711278
rect 390022 711042 390204 711278
rect 389604 710958 390204 711042
rect 389604 710722 389786 710958
rect 390022 710722 390204 710958
rect 386004 709438 386604 709460
rect 386004 709202 386186 709438
rect 386422 709202 386604 709438
rect 386004 709118 386604 709202
rect 386004 708882 386186 709118
rect 386422 708882 386604 709118
rect 382404 707598 383004 707620
rect 382404 707362 382586 707598
rect 382822 707362 383004 707598
rect 382404 707278 383004 707362
rect 382404 707042 382586 707278
rect 382822 707042 383004 707278
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 625254 372204 660698
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 589254 372204 624698
rect 371604 589018 371786 589254
rect 372022 589018 372204 589254
rect 371604 588934 372204 589018
rect 371604 588698 371786 588934
rect 372022 588698 372204 588934
rect 371604 553254 372204 588698
rect 371604 553018 371786 553254
rect 372022 553018 372204 553254
rect 371604 552934 372204 553018
rect 371604 552698 371786 552934
rect 372022 552698 372204 552934
rect 371604 517254 372204 552698
rect 371604 517018 371786 517254
rect 372022 517018 372204 517254
rect 371604 516934 372204 517018
rect 371604 516698 371786 516934
rect 372022 516698 372204 516934
rect 371604 481254 372204 516698
rect 371604 481018 371786 481254
rect 372022 481018 372204 481254
rect 371604 480934 372204 481018
rect 371604 480698 371786 480934
rect 372022 480698 372204 480934
rect 371604 445254 372204 480698
rect 371604 445018 371786 445254
rect 372022 445018 372204 445254
rect 371604 444934 372204 445018
rect 371604 444698 371786 444934
rect 372022 444698 372204 444934
rect 371604 409254 372204 444698
rect 371604 409018 371786 409254
rect 372022 409018 372204 409254
rect 371604 408934 372204 409018
rect 371604 408698 371786 408934
rect 372022 408698 372204 408934
rect 371604 373254 372204 408698
rect 371604 373018 371786 373254
rect 372022 373018 372204 373254
rect 371604 372934 372204 373018
rect 371604 372698 371786 372934
rect 372022 372698 372204 372934
rect 371604 337254 372204 372698
rect 371604 337018 371786 337254
rect 372022 337018 372204 337254
rect 371604 336934 372204 337018
rect 371604 336698 371786 336934
rect 372022 336698 372204 336934
rect 371604 301254 372204 336698
rect 378804 705758 379404 705780
rect 378804 705522 378986 705758
rect 379222 705522 379404 705758
rect 378804 705438 379404 705522
rect 378804 705202 378986 705438
rect 379222 705202 379404 705438
rect 378804 668454 379404 705202
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 378804 560454 379404 595898
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 378804 524454 379404 559898
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 378804 488454 379404 523898
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 452454 379404 487898
rect 378804 452218 378986 452454
rect 379222 452218 379404 452454
rect 378804 452134 379404 452218
rect 378804 451898 378986 452134
rect 379222 451898 379404 452134
rect 378804 416454 379404 451898
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 380454 379404 415898
rect 378804 380218 378986 380454
rect 379222 380218 379404 380454
rect 378804 380134 379404 380218
rect 378804 379898 378986 380134
rect 379222 379898 379404 380134
rect 378804 344454 379404 379898
rect 378804 344218 378986 344454
rect 379222 344218 379404 344454
rect 378804 344134 379404 344218
rect 378804 343898 378986 344134
rect 379222 343898 379404 344134
rect 376707 310860 376773 310861
rect 376707 310796 376708 310860
rect 376772 310796 376773 310860
rect 376707 310795 376773 310796
rect 376710 310589 376770 310795
rect 376707 310588 376773 310589
rect 376707 310524 376708 310588
rect 376772 310524 376773 310588
rect 376707 310523 376773 310524
rect 371604 301018 371786 301254
rect 372022 301018 372204 301254
rect 371604 300934 372204 301018
rect 371604 300698 371786 300934
rect 372022 300698 372204 300934
rect 371604 265254 372204 300698
rect 371604 265018 371786 265254
rect 372022 265018 372204 265254
rect 371604 264934 372204 265018
rect 371604 264698 371786 264934
rect 372022 264698 372204 264934
rect 371604 229254 372204 264698
rect 378804 308454 379404 343898
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 272454 379404 307898
rect 378804 272218 378986 272454
rect 379222 272218 379404 272454
rect 378804 272134 379404 272218
rect 378804 271898 378986 272134
rect 379222 271898 379404 272134
rect 376707 263940 376773 263941
rect 376707 263876 376708 263940
rect 376772 263876 376773 263940
rect 376707 263875 376773 263876
rect 376710 263669 376770 263875
rect 376707 263668 376773 263669
rect 376707 263604 376708 263668
rect 376772 263604 376773 263668
rect 376707 263603 376773 263604
rect 371604 229018 371786 229254
rect 372022 229018 372204 229254
rect 371604 228934 372204 229018
rect 371604 228698 371786 228934
rect 372022 228698 372204 228934
rect 371604 193254 372204 228698
rect 378804 236454 379404 271898
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 376707 217020 376773 217021
rect 376707 216956 376708 217020
rect 376772 216956 376773 217020
rect 376707 216955 376773 216956
rect 376710 216749 376770 216955
rect 376707 216748 376773 216749
rect 376707 216684 376708 216748
rect 376772 216684 376773 216748
rect 376707 216683 376773 216684
rect 371604 193018 371786 193254
rect 372022 193018 372204 193254
rect 371604 192934 372204 193018
rect 371604 192698 371786 192934
rect 372022 192698 372204 192934
rect 371604 157254 372204 192698
rect 378804 200454 379404 235898
rect 378804 200218 378986 200454
rect 379222 200218 379404 200454
rect 378804 200134 379404 200218
rect 378804 199898 378986 200134
rect 379222 199898 379404 200134
rect 376707 170100 376773 170101
rect 376707 170036 376708 170100
rect 376772 170036 376773 170100
rect 376707 170035 376773 170036
rect 376710 169829 376770 170035
rect 376707 169828 376773 169829
rect 376707 169764 376708 169828
rect 376772 169764 376773 169828
rect 376707 169763 376773 169764
rect 371604 157018 371786 157254
rect 372022 157018 372204 157254
rect 371604 156934 372204 157018
rect 371604 156698 371786 156934
rect 372022 156698 372204 156934
rect 371604 121254 372204 156698
rect 371604 121018 371786 121254
rect 372022 121018 372204 121254
rect 371604 120934 372204 121018
rect 371604 120698 371786 120934
rect 372022 120698 372204 120934
rect 371604 85254 372204 120698
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 378804 164454 379404 199898
rect 378804 164218 378986 164454
rect 379222 164218 379404 164454
rect 378804 164134 379404 164218
rect 378804 163898 378986 164134
rect 379222 163898 379404 164134
rect 378804 128454 379404 163898
rect 378804 128218 378986 128454
rect 379222 128218 379404 128454
rect 378804 128134 379404 128218
rect 378804 127898 378986 128134
rect 379222 127898 379404 128134
rect 378804 92454 379404 127898
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 376707 63884 376773 63885
rect 376707 63820 376708 63884
rect 376772 63820 376773 63884
rect 376707 63819 376773 63820
rect 376710 63613 376770 63819
rect 376707 63612 376773 63613
rect 376707 63548 376708 63612
rect 376772 63548 376773 63612
rect 376707 63547 376773 63548
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 376707 40356 376773 40357
rect 376707 40292 376708 40356
rect 376772 40292 376773 40356
rect 376707 40291 376773 40292
rect 376710 40085 376770 40291
rect 376707 40084 376773 40085
rect 376707 40020 376708 40084
rect 376772 40020 376773 40084
rect 376707 40019 376773 40020
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7022 353786 -6786
rect 354022 -7022 354204 -6786
rect 353604 -7106 354204 -7022
rect 353604 -7342 353786 -7106
rect 354022 -7342 354204 -7106
rect 353604 -7364 354204 -7342
rect 371604 -5866 372204 12698
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1266 379404 19898
rect 378804 -1502 378986 -1266
rect 379222 -1502 379404 -1266
rect 378804 -1586 379404 -1502
rect 378804 -1822 378986 -1586
rect 379222 -1822 379404 -1586
rect 378804 -1844 379404 -1822
rect 382404 672054 383004 707042
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 600054 383004 635498
rect 382404 599818 382586 600054
rect 382822 599818 383004 600054
rect 382404 599734 383004 599818
rect 382404 599498 382586 599734
rect 382822 599498 383004 599734
rect 382404 564054 383004 599498
rect 382404 563818 382586 564054
rect 382822 563818 383004 564054
rect 382404 563734 383004 563818
rect 382404 563498 382586 563734
rect 382822 563498 383004 563734
rect 382404 528054 383004 563498
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 382404 492054 383004 527498
rect 382404 491818 382586 492054
rect 382822 491818 383004 492054
rect 382404 491734 383004 491818
rect 382404 491498 382586 491734
rect 382822 491498 383004 491734
rect 382404 456054 383004 491498
rect 382404 455818 382586 456054
rect 382822 455818 383004 456054
rect 382404 455734 383004 455818
rect 382404 455498 382586 455734
rect 382822 455498 383004 455734
rect 382404 420054 383004 455498
rect 382404 419818 382586 420054
rect 382822 419818 383004 420054
rect 382404 419734 383004 419818
rect 382404 419498 382586 419734
rect 382822 419498 383004 419734
rect 382404 384054 383004 419498
rect 382404 383818 382586 384054
rect 382822 383818 383004 384054
rect 382404 383734 383004 383818
rect 382404 383498 382586 383734
rect 382822 383498 383004 383734
rect 382404 348054 383004 383498
rect 382404 347818 382586 348054
rect 382822 347818 383004 348054
rect 382404 347734 383004 347818
rect 382404 347498 382586 347734
rect 382822 347498 383004 347734
rect 382404 312054 383004 347498
rect 382404 311818 382586 312054
rect 382822 311818 383004 312054
rect 382404 311734 383004 311818
rect 382404 311498 382586 311734
rect 382822 311498 383004 311734
rect 382404 276054 383004 311498
rect 382404 275818 382586 276054
rect 382822 275818 383004 276054
rect 382404 275734 383004 275818
rect 382404 275498 382586 275734
rect 382822 275498 383004 275734
rect 382404 240054 383004 275498
rect 382404 239818 382586 240054
rect 382822 239818 383004 240054
rect 382404 239734 383004 239818
rect 382404 239498 382586 239734
rect 382822 239498 383004 239734
rect 382404 204054 383004 239498
rect 382404 203818 382586 204054
rect 382822 203818 383004 204054
rect 382404 203734 383004 203818
rect 382404 203498 382586 203734
rect 382822 203498 383004 203734
rect 382404 168054 383004 203498
rect 382404 167818 382586 168054
rect 382822 167818 383004 168054
rect 382404 167734 383004 167818
rect 382404 167498 382586 167734
rect 382822 167498 383004 167734
rect 382404 132054 383004 167498
rect 382404 131818 382586 132054
rect 382822 131818 383004 132054
rect 382404 131734 383004 131818
rect 382404 131498 382586 131734
rect 382822 131498 383004 131734
rect 382404 96054 383004 131498
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3106 383004 23498
rect 382404 -3342 382586 -3106
rect 382822 -3342 383004 -3106
rect 382404 -3426 383004 -3342
rect 382404 -3662 382586 -3426
rect 382822 -3662 383004 -3426
rect 382404 -3684 383004 -3662
rect 386004 675654 386604 708882
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 639654 386604 675098
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 386004 603654 386604 639098
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 567654 386604 603098
rect 386004 567418 386186 567654
rect 386422 567418 386604 567654
rect 386004 567334 386604 567418
rect 386004 567098 386186 567334
rect 386422 567098 386604 567334
rect 386004 531654 386604 567098
rect 386004 531418 386186 531654
rect 386422 531418 386604 531654
rect 386004 531334 386604 531418
rect 386004 531098 386186 531334
rect 386422 531098 386604 531334
rect 386004 495654 386604 531098
rect 386004 495418 386186 495654
rect 386422 495418 386604 495654
rect 386004 495334 386604 495418
rect 386004 495098 386186 495334
rect 386422 495098 386604 495334
rect 386004 459654 386604 495098
rect 386004 459418 386186 459654
rect 386422 459418 386604 459654
rect 386004 459334 386604 459418
rect 386004 459098 386186 459334
rect 386422 459098 386604 459334
rect 386004 423654 386604 459098
rect 386004 423418 386186 423654
rect 386422 423418 386604 423654
rect 386004 423334 386604 423418
rect 386004 423098 386186 423334
rect 386422 423098 386604 423334
rect 386004 387654 386604 423098
rect 386004 387418 386186 387654
rect 386422 387418 386604 387654
rect 386004 387334 386604 387418
rect 386004 387098 386186 387334
rect 386422 387098 386604 387334
rect 386004 351654 386604 387098
rect 386004 351418 386186 351654
rect 386422 351418 386604 351654
rect 386004 351334 386604 351418
rect 386004 351098 386186 351334
rect 386422 351098 386604 351334
rect 386004 315654 386604 351098
rect 386004 315418 386186 315654
rect 386422 315418 386604 315654
rect 386004 315334 386604 315418
rect 386004 315098 386186 315334
rect 386422 315098 386604 315334
rect 386004 279654 386604 315098
rect 386004 279418 386186 279654
rect 386422 279418 386604 279654
rect 386004 279334 386604 279418
rect 386004 279098 386186 279334
rect 386422 279098 386604 279334
rect 386004 243654 386604 279098
rect 386004 243418 386186 243654
rect 386422 243418 386604 243654
rect 386004 243334 386604 243418
rect 386004 243098 386186 243334
rect 386422 243098 386604 243334
rect 386004 207654 386604 243098
rect 386004 207418 386186 207654
rect 386422 207418 386604 207654
rect 386004 207334 386604 207418
rect 386004 207098 386186 207334
rect 386422 207098 386604 207334
rect 386004 171654 386604 207098
rect 386004 171418 386186 171654
rect 386422 171418 386604 171654
rect 386004 171334 386604 171418
rect 386004 171098 386186 171334
rect 386422 171098 386604 171334
rect 386004 135654 386604 171098
rect 386004 135418 386186 135654
rect 386422 135418 386604 135654
rect 386004 135334 386604 135418
rect 386004 135098 386186 135334
rect 386422 135098 386604 135334
rect 386004 99654 386604 135098
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -4946 386604 27098
rect 386004 -5182 386186 -4946
rect 386422 -5182 386604 -4946
rect 386004 -5266 386604 -5182
rect 386004 -5502 386186 -5266
rect 386422 -5502 386604 -5266
rect 386004 -5524 386604 -5502
rect 389604 679254 390204 710722
rect 407604 710358 408204 711300
rect 407604 710122 407786 710358
rect 408022 710122 408204 710358
rect 407604 710038 408204 710122
rect 407604 709802 407786 710038
rect 408022 709802 408204 710038
rect 404004 708518 404604 709460
rect 404004 708282 404186 708518
rect 404422 708282 404604 708518
rect 404004 708198 404604 708282
rect 404004 707962 404186 708198
rect 404422 707962 404604 708198
rect 400404 706678 401004 707620
rect 400404 706442 400586 706678
rect 400822 706442 401004 706678
rect 400404 706358 401004 706442
rect 400404 706122 400586 706358
rect 400822 706122 401004 706358
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 389604 607254 390204 642698
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 389604 571254 390204 606698
rect 389604 571018 389786 571254
rect 390022 571018 390204 571254
rect 389604 570934 390204 571018
rect 389604 570698 389786 570934
rect 390022 570698 390204 570934
rect 389604 535254 390204 570698
rect 389604 535018 389786 535254
rect 390022 535018 390204 535254
rect 389604 534934 390204 535018
rect 389604 534698 389786 534934
rect 390022 534698 390204 534934
rect 389604 499254 390204 534698
rect 389604 499018 389786 499254
rect 390022 499018 390204 499254
rect 389604 498934 390204 499018
rect 389604 498698 389786 498934
rect 390022 498698 390204 498934
rect 389604 463254 390204 498698
rect 389604 463018 389786 463254
rect 390022 463018 390204 463254
rect 389604 462934 390204 463018
rect 389604 462698 389786 462934
rect 390022 462698 390204 462934
rect 389604 427254 390204 462698
rect 389604 427018 389786 427254
rect 390022 427018 390204 427254
rect 389604 426934 390204 427018
rect 389604 426698 389786 426934
rect 390022 426698 390204 426934
rect 389604 391254 390204 426698
rect 389604 391018 389786 391254
rect 390022 391018 390204 391254
rect 389604 390934 390204 391018
rect 389604 390698 389786 390934
rect 390022 390698 390204 390934
rect 389604 355254 390204 390698
rect 389604 355018 389786 355254
rect 390022 355018 390204 355254
rect 389604 354934 390204 355018
rect 389604 354698 389786 354934
rect 390022 354698 390204 354934
rect 389604 319254 390204 354698
rect 389604 319018 389786 319254
rect 390022 319018 390204 319254
rect 389604 318934 390204 319018
rect 389604 318698 389786 318934
rect 390022 318698 390204 318934
rect 389604 283254 390204 318698
rect 389604 283018 389786 283254
rect 390022 283018 390204 283254
rect 389604 282934 390204 283018
rect 389604 282698 389786 282934
rect 390022 282698 390204 282934
rect 389604 247254 390204 282698
rect 389604 247018 389786 247254
rect 390022 247018 390204 247254
rect 389604 246934 390204 247018
rect 389604 246698 389786 246934
rect 390022 246698 390204 246934
rect 389604 211254 390204 246698
rect 389604 211018 389786 211254
rect 390022 211018 390204 211254
rect 389604 210934 390204 211018
rect 389604 210698 389786 210934
rect 390022 210698 390204 210934
rect 389604 175254 390204 210698
rect 389604 175018 389786 175254
rect 390022 175018 390204 175254
rect 389604 174934 390204 175018
rect 389604 174698 389786 174934
rect 390022 174698 390204 174934
rect 389604 139254 390204 174698
rect 389604 139018 389786 139254
rect 390022 139018 390204 139254
rect 389604 138934 390204 139018
rect 389604 138698 389786 138934
rect 390022 138698 390204 138934
rect 389604 103254 390204 138698
rect 389604 103018 389786 103254
rect 390022 103018 390204 103254
rect 389604 102934 390204 103018
rect 389604 102698 389786 102934
rect 390022 102698 390204 102934
rect 389604 67254 390204 102698
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6102 371786 -5866
rect 372022 -6102 372204 -5866
rect 371604 -6186 372204 -6102
rect 371604 -6422 371786 -6186
rect 372022 -6422 372204 -6186
rect 371604 -7364 372204 -6422
rect 389604 -6786 390204 30698
rect 396804 704838 397404 705780
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 396804 470454 397404 505898
rect 396804 470218 396986 470454
rect 397222 470218 397404 470454
rect 396804 470134 397404 470218
rect 396804 469898 396986 470134
rect 397222 469898 397404 470134
rect 396804 434454 397404 469898
rect 396804 434218 396986 434454
rect 397222 434218 397404 434454
rect 396804 434134 397404 434218
rect 396804 433898 396986 434134
rect 397222 433898 397404 434134
rect 396804 398454 397404 433898
rect 396804 398218 396986 398454
rect 397222 398218 397404 398454
rect 396804 398134 397404 398218
rect 396804 397898 396986 398134
rect 397222 397898 397404 398134
rect 396804 362454 397404 397898
rect 396804 362218 396986 362454
rect 397222 362218 397404 362454
rect 396804 362134 397404 362218
rect 396804 361898 396986 362134
rect 397222 361898 397404 362134
rect 396804 326454 397404 361898
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 396804 290454 397404 325898
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 396804 254454 397404 289898
rect 396804 254218 396986 254454
rect 397222 254218 397404 254454
rect 396804 254134 397404 254218
rect 396804 253898 396986 254134
rect 397222 253898 397404 254134
rect 396804 218454 397404 253898
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 182454 397404 217898
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1844 397404 -902
rect 400404 690054 401004 706122
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 510054 401004 545498
rect 400404 509818 400586 510054
rect 400822 509818 401004 510054
rect 400404 509734 401004 509818
rect 400404 509498 400586 509734
rect 400822 509498 401004 509734
rect 400404 474054 401004 509498
rect 400404 473818 400586 474054
rect 400822 473818 401004 474054
rect 400404 473734 401004 473818
rect 400404 473498 400586 473734
rect 400822 473498 401004 473734
rect 400404 438054 401004 473498
rect 400404 437818 400586 438054
rect 400822 437818 401004 438054
rect 400404 437734 401004 437818
rect 400404 437498 400586 437734
rect 400822 437498 401004 437734
rect 400404 402054 401004 437498
rect 400404 401818 400586 402054
rect 400822 401818 401004 402054
rect 400404 401734 401004 401818
rect 400404 401498 400586 401734
rect 400822 401498 401004 401734
rect 400404 366054 401004 401498
rect 400404 365818 400586 366054
rect 400822 365818 401004 366054
rect 400404 365734 401004 365818
rect 400404 365498 400586 365734
rect 400822 365498 401004 365734
rect 400404 330054 401004 365498
rect 400404 329818 400586 330054
rect 400822 329818 401004 330054
rect 400404 329734 401004 329818
rect 400404 329498 400586 329734
rect 400822 329498 401004 329734
rect 400404 294054 401004 329498
rect 400404 293818 400586 294054
rect 400822 293818 401004 294054
rect 400404 293734 401004 293818
rect 400404 293498 400586 293734
rect 400822 293498 401004 293734
rect 400404 258054 401004 293498
rect 400404 257818 400586 258054
rect 400822 257818 401004 258054
rect 400404 257734 401004 257818
rect 400404 257498 400586 257734
rect 400822 257498 401004 257734
rect 400404 222054 401004 257498
rect 400404 221818 400586 222054
rect 400822 221818 401004 222054
rect 400404 221734 401004 221818
rect 400404 221498 400586 221734
rect 400822 221498 401004 221734
rect 400404 186054 401004 221498
rect 400404 185818 400586 186054
rect 400822 185818 401004 186054
rect 400404 185734 401004 185818
rect 400404 185498 400586 185734
rect 400822 185498 401004 185734
rect 400404 150054 401004 185498
rect 400404 149818 400586 150054
rect 400822 149818 401004 150054
rect 400404 149734 401004 149818
rect 400404 149498 400586 149734
rect 400822 149498 401004 149734
rect 400404 114054 401004 149498
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2186 401004 5498
rect 400404 -2422 400586 -2186
rect 400822 -2422 401004 -2186
rect 400404 -2506 401004 -2422
rect 400404 -2742 400586 -2506
rect 400822 -2742 401004 -2506
rect 400404 -3684 401004 -2742
rect 404004 693654 404604 707962
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 513654 404604 549098
rect 404004 513418 404186 513654
rect 404422 513418 404604 513654
rect 404004 513334 404604 513418
rect 404004 513098 404186 513334
rect 404422 513098 404604 513334
rect 404004 477654 404604 513098
rect 404004 477418 404186 477654
rect 404422 477418 404604 477654
rect 404004 477334 404604 477418
rect 404004 477098 404186 477334
rect 404422 477098 404604 477334
rect 404004 441654 404604 477098
rect 404004 441418 404186 441654
rect 404422 441418 404604 441654
rect 404004 441334 404604 441418
rect 404004 441098 404186 441334
rect 404422 441098 404604 441334
rect 404004 405654 404604 441098
rect 404004 405418 404186 405654
rect 404422 405418 404604 405654
rect 404004 405334 404604 405418
rect 404004 405098 404186 405334
rect 404422 405098 404604 405334
rect 404004 369654 404604 405098
rect 404004 369418 404186 369654
rect 404422 369418 404604 369654
rect 404004 369334 404604 369418
rect 404004 369098 404186 369334
rect 404422 369098 404604 369334
rect 404004 333654 404604 369098
rect 404004 333418 404186 333654
rect 404422 333418 404604 333654
rect 404004 333334 404604 333418
rect 404004 333098 404186 333334
rect 404422 333098 404604 333334
rect 404004 297654 404604 333098
rect 404004 297418 404186 297654
rect 404422 297418 404604 297654
rect 404004 297334 404604 297418
rect 404004 297098 404186 297334
rect 404422 297098 404604 297334
rect 404004 261654 404604 297098
rect 404004 261418 404186 261654
rect 404422 261418 404604 261654
rect 404004 261334 404604 261418
rect 404004 261098 404186 261334
rect 404422 261098 404604 261334
rect 404004 225654 404604 261098
rect 404004 225418 404186 225654
rect 404422 225418 404604 225654
rect 404004 225334 404604 225418
rect 404004 225098 404186 225334
rect 404422 225098 404604 225334
rect 404004 189654 404604 225098
rect 404004 189418 404186 189654
rect 404422 189418 404604 189654
rect 404004 189334 404604 189418
rect 404004 189098 404186 189334
rect 404422 189098 404604 189334
rect 404004 153654 404604 189098
rect 404004 153418 404186 153654
rect 404422 153418 404604 153654
rect 404004 153334 404604 153418
rect 404004 153098 404186 153334
rect 404422 153098 404604 153334
rect 404004 117654 404604 153098
rect 404004 117418 404186 117654
rect 404422 117418 404604 117654
rect 404004 117334 404604 117418
rect 404004 117098 404186 117334
rect 404422 117098 404604 117334
rect 404004 81654 404604 117098
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4026 404604 9098
rect 404004 -4262 404186 -4026
rect 404422 -4262 404604 -4026
rect 404004 -4346 404604 -4262
rect 404004 -4582 404186 -4346
rect 404422 -4582 404604 -4346
rect 404004 -5524 404604 -4582
rect 407604 697254 408204 709802
rect 425604 711278 426204 711300
rect 425604 711042 425786 711278
rect 426022 711042 426204 711278
rect 425604 710958 426204 711042
rect 425604 710722 425786 710958
rect 426022 710722 426204 710958
rect 422004 709438 422604 709460
rect 422004 709202 422186 709438
rect 422422 709202 422604 709438
rect 422004 709118 422604 709202
rect 422004 708882 422186 709118
rect 422422 708882 422604 709118
rect 418404 707598 419004 707620
rect 418404 707362 418586 707598
rect 418822 707362 419004 707598
rect 418404 707278 419004 707362
rect 418404 707042 418586 707278
rect 418822 707042 419004 707278
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 553254 408204 588698
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 517254 408204 552698
rect 407604 517018 407786 517254
rect 408022 517018 408204 517254
rect 407604 516934 408204 517018
rect 407604 516698 407786 516934
rect 408022 516698 408204 516934
rect 407604 481254 408204 516698
rect 407604 481018 407786 481254
rect 408022 481018 408204 481254
rect 407604 480934 408204 481018
rect 407604 480698 407786 480934
rect 408022 480698 408204 480934
rect 407604 445254 408204 480698
rect 407604 445018 407786 445254
rect 408022 445018 408204 445254
rect 407604 444934 408204 445018
rect 407604 444698 407786 444934
rect 408022 444698 408204 444934
rect 407604 409254 408204 444698
rect 407604 409018 407786 409254
rect 408022 409018 408204 409254
rect 407604 408934 408204 409018
rect 407604 408698 407786 408934
rect 408022 408698 408204 408934
rect 407604 373254 408204 408698
rect 407604 373018 407786 373254
rect 408022 373018 408204 373254
rect 407604 372934 408204 373018
rect 407604 372698 407786 372934
rect 408022 372698 408204 372934
rect 407604 337254 408204 372698
rect 407604 337018 407786 337254
rect 408022 337018 408204 337254
rect 407604 336934 408204 337018
rect 407604 336698 407786 336934
rect 408022 336698 408204 336934
rect 407604 301254 408204 336698
rect 407604 301018 407786 301254
rect 408022 301018 408204 301254
rect 407604 300934 408204 301018
rect 407604 300698 407786 300934
rect 408022 300698 408204 300934
rect 407604 265254 408204 300698
rect 407604 265018 407786 265254
rect 408022 265018 408204 265254
rect 407604 264934 408204 265018
rect 407604 264698 407786 264934
rect 408022 264698 408204 264934
rect 407604 229254 408204 264698
rect 407604 229018 407786 229254
rect 408022 229018 408204 229254
rect 407604 228934 408204 229018
rect 407604 228698 407786 228934
rect 408022 228698 408204 228934
rect 407604 193254 408204 228698
rect 407604 193018 407786 193254
rect 408022 193018 408204 193254
rect 407604 192934 408204 193018
rect 407604 192698 407786 192934
rect 408022 192698 408204 192934
rect 407604 157254 408204 192698
rect 407604 157018 407786 157254
rect 408022 157018 408204 157254
rect 407604 156934 408204 157018
rect 407604 156698 407786 156934
rect 408022 156698 408204 156934
rect 407604 121254 408204 156698
rect 407604 121018 407786 121254
rect 408022 121018 408204 121254
rect 407604 120934 408204 121018
rect 407604 120698 407786 120934
rect 408022 120698 408204 120934
rect 407604 85254 408204 120698
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7022 389786 -6786
rect 390022 -7022 390204 -6786
rect 389604 -7106 390204 -7022
rect 389604 -7342 389786 -7106
rect 390022 -7342 390204 -7106
rect 389604 -7364 390204 -7342
rect 407604 -5866 408204 12698
rect 414804 705758 415404 705780
rect 414804 705522 414986 705758
rect 415222 705522 415404 705758
rect 414804 705438 415404 705522
rect 414804 705202 414986 705438
rect 415222 705202 415404 705438
rect 414804 668454 415404 705202
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 380454 415404 415898
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 272454 415404 307898
rect 414804 272218 414986 272454
rect 415222 272218 415404 272454
rect 414804 272134 415404 272218
rect 414804 271898 414986 272134
rect 415222 271898 415404 272134
rect 414804 236454 415404 271898
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1266 415404 19898
rect 414804 -1502 414986 -1266
rect 415222 -1502 415404 -1266
rect 414804 -1586 415404 -1502
rect 414804 -1822 414986 -1586
rect 415222 -1822 415404 -1586
rect 414804 -1844 415404 -1822
rect 418404 672054 419004 707042
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 528054 419004 563498
rect 418404 527818 418586 528054
rect 418822 527818 419004 528054
rect 418404 527734 419004 527818
rect 418404 527498 418586 527734
rect 418822 527498 419004 527734
rect 418404 492054 419004 527498
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 456054 419004 491498
rect 418404 455818 418586 456054
rect 418822 455818 419004 456054
rect 418404 455734 419004 455818
rect 418404 455498 418586 455734
rect 418822 455498 419004 455734
rect 418404 420054 419004 455498
rect 418404 419818 418586 420054
rect 418822 419818 419004 420054
rect 418404 419734 419004 419818
rect 418404 419498 418586 419734
rect 418822 419498 419004 419734
rect 418404 384054 419004 419498
rect 418404 383818 418586 384054
rect 418822 383818 419004 384054
rect 418404 383734 419004 383818
rect 418404 383498 418586 383734
rect 418822 383498 419004 383734
rect 418404 348054 419004 383498
rect 418404 347818 418586 348054
rect 418822 347818 419004 348054
rect 418404 347734 419004 347818
rect 418404 347498 418586 347734
rect 418822 347498 419004 347734
rect 418404 312054 419004 347498
rect 418404 311818 418586 312054
rect 418822 311818 419004 312054
rect 418404 311734 419004 311818
rect 418404 311498 418586 311734
rect 418822 311498 419004 311734
rect 418404 276054 419004 311498
rect 418404 275818 418586 276054
rect 418822 275818 419004 276054
rect 418404 275734 419004 275818
rect 418404 275498 418586 275734
rect 418822 275498 419004 275734
rect 418404 240054 419004 275498
rect 418404 239818 418586 240054
rect 418822 239818 419004 240054
rect 418404 239734 419004 239818
rect 418404 239498 418586 239734
rect 418822 239498 419004 239734
rect 418404 204054 419004 239498
rect 418404 203818 418586 204054
rect 418822 203818 419004 204054
rect 418404 203734 419004 203818
rect 418404 203498 418586 203734
rect 418822 203498 419004 203734
rect 418404 168054 419004 203498
rect 418404 167818 418586 168054
rect 418822 167818 419004 168054
rect 418404 167734 419004 167818
rect 418404 167498 418586 167734
rect 418822 167498 419004 167734
rect 418404 132054 419004 167498
rect 418404 131818 418586 132054
rect 418822 131818 419004 132054
rect 418404 131734 419004 131818
rect 418404 131498 418586 131734
rect 418822 131498 419004 131734
rect 418404 96054 419004 131498
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3106 419004 23498
rect 418404 -3342 418586 -3106
rect 418822 -3342 419004 -3106
rect 418404 -3426 419004 -3342
rect 418404 -3662 418586 -3426
rect 418822 -3662 419004 -3426
rect 418404 -3684 419004 -3662
rect 422004 675654 422604 708882
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 567654 422604 603098
rect 422004 567418 422186 567654
rect 422422 567418 422604 567654
rect 422004 567334 422604 567418
rect 422004 567098 422186 567334
rect 422422 567098 422604 567334
rect 422004 531654 422604 567098
rect 422004 531418 422186 531654
rect 422422 531418 422604 531654
rect 422004 531334 422604 531418
rect 422004 531098 422186 531334
rect 422422 531098 422604 531334
rect 422004 495654 422604 531098
rect 422004 495418 422186 495654
rect 422422 495418 422604 495654
rect 422004 495334 422604 495418
rect 422004 495098 422186 495334
rect 422422 495098 422604 495334
rect 422004 459654 422604 495098
rect 422004 459418 422186 459654
rect 422422 459418 422604 459654
rect 422004 459334 422604 459418
rect 422004 459098 422186 459334
rect 422422 459098 422604 459334
rect 422004 423654 422604 459098
rect 422004 423418 422186 423654
rect 422422 423418 422604 423654
rect 422004 423334 422604 423418
rect 422004 423098 422186 423334
rect 422422 423098 422604 423334
rect 422004 387654 422604 423098
rect 422004 387418 422186 387654
rect 422422 387418 422604 387654
rect 422004 387334 422604 387418
rect 422004 387098 422186 387334
rect 422422 387098 422604 387334
rect 422004 351654 422604 387098
rect 422004 351418 422186 351654
rect 422422 351418 422604 351654
rect 422004 351334 422604 351418
rect 422004 351098 422186 351334
rect 422422 351098 422604 351334
rect 422004 315654 422604 351098
rect 422004 315418 422186 315654
rect 422422 315418 422604 315654
rect 422004 315334 422604 315418
rect 422004 315098 422186 315334
rect 422422 315098 422604 315334
rect 422004 279654 422604 315098
rect 422004 279418 422186 279654
rect 422422 279418 422604 279654
rect 422004 279334 422604 279418
rect 422004 279098 422186 279334
rect 422422 279098 422604 279334
rect 422004 243654 422604 279098
rect 422004 243418 422186 243654
rect 422422 243418 422604 243654
rect 422004 243334 422604 243418
rect 422004 243098 422186 243334
rect 422422 243098 422604 243334
rect 422004 207654 422604 243098
rect 422004 207418 422186 207654
rect 422422 207418 422604 207654
rect 422004 207334 422604 207418
rect 422004 207098 422186 207334
rect 422422 207098 422604 207334
rect 422004 171654 422604 207098
rect 422004 171418 422186 171654
rect 422422 171418 422604 171654
rect 422004 171334 422604 171418
rect 422004 171098 422186 171334
rect 422422 171098 422604 171334
rect 422004 135654 422604 171098
rect 422004 135418 422186 135654
rect 422422 135418 422604 135654
rect 422004 135334 422604 135418
rect 422004 135098 422186 135334
rect 422422 135098 422604 135334
rect 422004 99654 422604 135098
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -4946 422604 27098
rect 422004 -5182 422186 -4946
rect 422422 -5182 422604 -4946
rect 422004 -5266 422604 -5182
rect 422004 -5502 422186 -5266
rect 422422 -5502 422604 -5266
rect 422004 -5524 422604 -5502
rect 425604 679254 426204 710722
rect 443604 710358 444204 711300
rect 443604 710122 443786 710358
rect 444022 710122 444204 710358
rect 443604 710038 444204 710122
rect 443604 709802 443786 710038
rect 444022 709802 444204 710038
rect 440004 708518 440604 709460
rect 440004 708282 440186 708518
rect 440422 708282 440604 708518
rect 440004 708198 440604 708282
rect 440004 707962 440186 708198
rect 440422 707962 440604 708198
rect 436404 706678 437004 707620
rect 436404 706442 436586 706678
rect 436822 706442 437004 706678
rect 436404 706358 437004 706442
rect 436404 706122 436586 706358
rect 436822 706122 437004 706358
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 571254 426204 606698
rect 425604 571018 425786 571254
rect 426022 571018 426204 571254
rect 425604 570934 426204 571018
rect 425604 570698 425786 570934
rect 426022 570698 426204 570934
rect 425604 535254 426204 570698
rect 425604 535018 425786 535254
rect 426022 535018 426204 535254
rect 425604 534934 426204 535018
rect 425604 534698 425786 534934
rect 426022 534698 426204 534934
rect 425604 499254 426204 534698
rect 425604 499018 425786 499254
rect 426022 499018 426204 499254
rect 425604 498934 426204 499018
rect 425604 498698 425786 498934
rect 426022 498698 426204 498934
rect 425604 463254 426204 498698
rect 425604 463018 425786 463254
rect 426022 463018 426204 463254
rect 425604 462934 426204 463018
rect 425604 462698 425786 462934
rect 426022 462698 426204 462934
rect 425604 427254 426204 462698
rect 425604 427018 425786 427254
rect 426022 427018 426204 427254
rect 425604 426934 426204 427018
rect 425604 426698 425786 426934
rect 426022 426698 426204 426934
rect 425604 391254 426204 426698
rect 425604 391018 425786 391254
rect 426022 391018 426204 391254
rect 425604 390934 426204 391018
rect 425604 390698 425786 390934
rect 426022 390698 426204 390934
rect 425604 355254 426204 390698
rect 425604 355018 425786 355254
rect 426022 355018 426204 355254
rect 425604 354934 426204 355018
rect 425604 354698 425786 354934
rect 426022 354698 426204 354934
rect 425604 319254 426204 354698
rect 425604 319018 425786 319254
rect 426022 319018 426204 319254
rect 425604 318934 426204 319018
rect 425604 318698 425786 318934
rect 426022 318698 426204 318934
rect 425604 283254 426204 318698
rect 425604 283018 425786 283254
rect 426022 283018 426204 283254
rect 425604 282934 426204 283018
rect 425604 282698 425786 282934
rect 426022 282698 426204 282934
rect 425604 247254 426204 282698
rect 425604 247018 425786 247254
rect 426022 247018 426204 247254
rect 425604 246934 426204 247018
rect 425604 246698 425786 246934
rect 426022 246698 426204 246934
rect 425604 211254 426204 246698
rect 425604 211018 425786 211254
rect 426022 211018 426204 211254
rect 425604 210934 426204 211018
rect 425604 210698 425786 210934
rect 426022 210698 426204 210934
rect 425604 175254 426204 210698
rect 425604 175018 425786 175254
rect 426022 175018 426204 175254
rect 425604 174934 426204 175018
rect 425604 174698 425786 174934
rect 426022 174698 426204 174934
rect 425604 139254 426204 174698
rect 425604 139018 425786 139254
rect 426022 139018 426204 139254
rect 425604 138934 426204 139018
rect 425604 138698 425786 138934
rect 426022 138698 426204 138934
rect 425604 103254 426204 138698
rect 425604 103018 425786 103254
rect 426022 103018 426204 103254
rect 425604 102934 426204 103018
rect 425604 102698 425786 102934
rect 426022 102698 426204 102934
rect 425604 67254 426204 102698
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6102 407786 -5866
rect 408022 -6102 408204 -5866
rect 407604 -6186 408204 -6102
rect 407604 -6422 407786 -6186
rect 408022 -6422 408204 -6186
rect 407604 -7364 408204 -6422
rect 425604 -6786 426204 30698
rect 432804 704838 433404 705780
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 506454 433404 541898
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 470454 433404 505898
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 254454 433404 289898
rect 432804 254218 432986 254454
rect 433222 254218 433404 254454
rect 432804 254134 433404 254218
rect 432804 253898 432986 254134
rect 433222 253898 433404 254134
rect 432804 218454 433404 253898
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 182454 433404 217898
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1844 433404 -902
rect 436404 690054 437004 706122
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 582054 437004 617498
rect 436404 581818 436586 582054
rect 436822 581818 437004 582054
rect 436404 581734 437004 581818
rect 436404 581498 436586 581734
rect 436822 581498 437004 581734
rect 436404 546054 437004 581498
rect 436404 545818 436586 546054
rect 436822 545818 437004 546054
rect 436404 545734 437004 545818
rect 436404 545498 436586 545734
rect 436822 545498 437004 545734
rect 436404 510054 437004 545498
rect 436404 509818 436586 510054
rect 436822 509818 437004 510054
rect 436404 509734 437004 509818
rect 436404 509498 436586 509734
rect 436822 509498 437004 509734
rect 436404 474054 437004 509498
rect 436404 473818 436586 474054
rect 436822 473818 437004 474054
rect 436404 473734 437004 473818
rect 436404 473498 436586 473734
rect 436822 473498 437004 473734
rect 436404 438054 437004 473498
rect 436404 437818 436586 438054
rect 436822 437818 437004 438054
rect 436404 437734 437004 437818
rect 436404 437498 436586 437734
rect 436822 437498 437004 437734
rect 436404 402054 437004 437498
rect 436404 401818 436586 402054
rect 436822 401818 437004 402054
rect 436404 401734 437004 401818
rect 436404 401498 436586 401734
rect 436822 401498 437004 401734
rect 436404 366054 437004 401498
rect 436404 365818 436586 366054
rect 436822 365818 437004 366054
rect 436404 365734 437004 365818
rect 436404 365498 436586 365734
rect 436822 365498 437004 365734
rect 436404 330054 437004 365498
rect 436404 329818 436586 330054
rect 436822 329818 437004 330054
rect 436404 329734 437004 329818
rect 436404 329498 436586 329734
rect 436822 329498 437004 329734
rect 436404 294054 437004 329498
rect 436404 293818 436586 294054
rect 436822 293818 437004 294054
rect 436404 293734 437004 293818
rect 436404 293498 436586 293734
rect 436822 293498 437004 293734
rect 436404 258054 437004 293498
rect 436404 257818 436586 258054
rect 436822 257818 437004 258054
rect 436404 257734 437004 257818
rect 436404 257498 436586 257734
rect 436822 257498 437004 257734
rect 436404 222054 437004 257498
rect 436404 221818 436586 222054
rect 436822 221818 437004 222054
rect 436404 221734 437004 221818
rect 436404 221498 436586 221734
rect 436822 221498 437004 221734
rect 436404 186054 437004 221498
rect 436404 185818 436586 186054
rect 436822 185818 437004 186054
rect 436404 185734 437004 185818
rect 436404 185498 436586 185734
rect 436822 185498 437004 185734
rect 436404 150054 437004 185498
rect 436404 149818 436586 150054
rect 436822 149818 437004 150054
rect 436404 149734 437004 149818
rect 436404 149498 436586 149734
rect 436822 149498 437004 149734
rect 436404 114054 437004 149498
rect 436404 113818 436586 114054
rect 436822 113818 437004 114054
rect 436404 113734 437004 113818
rect 436404 113498 436586 113734
rect 436822 113498 437004 113734
rect 436404 78054 437004 113498
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2186 437004 5498
rect 436404 -2422 436586 -2186
rect 436822 -2422 437004 -2186
rect 436404 -2506 437004 -2422
rect 436404 -2742 436586 -2506
rect 436822 -2742 437004 -2506
rect 436404 -3684 437004 -2742
rect 440004 693654 440604 707962
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 621654 440604 657098
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 585654 440604 621098
rect 440004 585418 440186 585654
rect 440422 585418 440604 585654
rect 440004 585334 440604 585418
rect 440004 585098 440186 585334
rect 440422 585098 440604 585334
rect 440004 549654 440604 585098
rect 440004 549418 440186 549654
rect 440422 549418 440604 549654
rect 440004 549334 440604 549418
rect 440004 549098 440186 549334
rect 440422 549098 440604 549334
rect 440004 513654 440604 549098
rect 440004 513418 440186 513654
rect 440422 513418 440604 513654
rect 440004 513334 440604 513418
rect 440004 513098 440186 513334
rect 440422 513098 440604 513334
rect 440004 477654 440604 513098
rect 440004 477418 440186 477654
rect 440422 477418 440604 477654
rect 440004 477334 440604 477418
rect 440004 477098 440186 477334
rect 440422 477098 440604 477334
rect 440004 441654 440604 477098
rect 440004 441418 440186 441654
rect 440422 441418 440604 441654
rect 440004 441334 440604 441418
rect 440004 441098 440186 441334
rect 440422 441098 440604 441334
rect 440004 405654 440604 441098
rect 440004 405418 440186 405654
rect 440422 405418 440604 405654
rect 440004 405334 440604 405418
rect 440004 405098 440186 405334
rect 440422 405098 440604 405334
rect 440004 369654 440604 405098
rect 440004 369418 440186 369654
rect 440422 369418 440604 369654
rect 440004 369334 440604 369418
rect 440004 369098 440186 369334
rect 440422 369098 440604 369334
rect 440004 333654 440604 369098
rect 440004 333418 440186 333654
rect 440422 333418 440604 333654
rect 440004 333334 440604 333418
rect 440004 333098 440186 333334
rect 440422 333098 440604 333334
rect 440004 297654 440604 333098
rect 440004 297418 440186 297654
rect 440422 297418 440604 297654
rect 440004 297334 440604 297418
rect 440004 297098 440186 297334
rect 440422 297098 440604 297334
rect 440004 261654 440604 297098
rect 440004 261418 440186 261654
rect 440422 261418 440604 261654
rect 440004 261334 440604 261418
rect 440004 261098 440186 261334
rect 440422 261098 440604 261334
rect 440004 225654 440604 261098
rect 440004 225418 440186 225654
rect 440422 225418 440604 225654
rect 440004 225334 440604 225418
rect 440004 225098 440186 225334
rect 440422 225098 440604 225334
rect 440004 189654 440604 225098
rect 440004 189418 440186 189654
rect 440422 189418 440604 189654
rect 440004 189334 440604 189418
rect 440004 189098 440186 189334
rect 440422 189098 440604 189334
rect 440004 153654 440604 189098
rect 440004 153418 440186 153654
rect 440422 153418 440604 153654
rect 440004 153334 440604 153418
rect 440004 153098 440186 153334
rect 440422 153098 440604 153334
rect 440004 117654 440604 153098
rect 440004 117418 440186 117654
rect 440422 117418 440604 117654
rect 440004 117334 440604 117418
rect 440004 117098 440186 117334
rect 440422 117098 440604 117334
rect 440004 81654 440604 117098
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4026 440604 9098
rect 440004 -4262 440186 -4026
rect 440422 -4262 440604 -4026
rect 440004 -4346 440604 -4262
rect 440004 -4582 440186 -4346
rect 440422 -4582 440604 -4346
rect 440004 -5524 440604 -4582
rect 443604 697254 444204 709802
rect 461604 711278 462204 711300
rect 461604 711042 461786 711278
rect 462022 711042 462204 711278
rect 461604 710958 462204 711042
rect 461604 710722 461786 710958
rect 462022 710722 462204 710958
rect 458004 709438 458604 709460
rect 458004 709202 458186 709438
rect 458422 709202 458604 709438
rect 458004 709118 458604 709202
rect 458004 708882 458186 709118
rect 458422 708882 458604 709118
rect 454404 707598 455004 707620
rect 454404 707362 454586 707598
rect 454822 707362 455004 707598
rect 454404 707278 455004 707362
rect 454404 707042 454586 707278
rect 454822 707042 455004 707278
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 589254 444204 624698
rect 443604 589018 443786 589254
rect 444022 589018 444204 589254
rect 443604 588934 444204 589018
rect 443604 588698 443786 588934
rect 444022 588698 444204 588934
rect 443604 553254 444204 588698
rect 443604 553018 443786 553254
rect 444022 553018 444204 553254
rect 443604 552934 444204 553018
rect 443604 552698 443786 552934
rect 444022 552698 444204 552934
rect 443604 517254 444204 552698
rect 443604 517018 443786 517254
rect 444022 517018 444204 517254
rect 443604 516934 444204 517018
rect 443604 516698 443786 516934
rect 444022 516698 444204 516934
rect 443604 481254 444204 516698
rect 443604 481018 443786 481254
rect 444022 481018 444204 481254
rect 443604 480934 444204 481018
rect 443604 480698 443786 480934
rect 444022 480698 444204 480934
rect 443604 445254 444204 480698
rect 443604 445018 443786 445254
rect 444022 445018 444204 445254
rect 443604 444934 444204 445018
rect 443604 444698 443786 444934
rect 444022 444698 444204 444934
rect 443604 409254 444204 444698
rect 443604 409018 443786 409254
rect 444022 409018 444204 409254
rect 443604 408934 444204 409018
rect 443604 408698 443786 408934
rect 444022 408698 444204 408934
rect 443604 373254 444204 408698
rect 443604 373018 443786 373254
rect 444022 373018 444204 373254
rect 443604 372934 444204 373018
rect 443604 372698 443786 372934
rect 444022 372698 444204 372934
rect 443604 337254 444204 372698
rect 443604 337018 443786 337254
rect 444022 337018 444204 337254
rect 443604 336934 444204 337018
rect 443604 336698 443786 336934
rect 444022 336698 444204 336934
rect 443604 301254 444204 336698
rect 443604 301018 443786 301254
rect 444022 301018 444204 301254
rect 443604 300934 444204 301018
rect 443604 300698 443786 300934
rect 444022 300698 444204 300934
rect 443604 265254 444204 300698
rect 443604 265018 443786 265254
rect 444022 265018 444204 265254
rect 443604 264934 444204 265018
rect 443604 264698 443786 264934
rect 444022 264698 444204 264934
rect 443604 229254 444204 264698
rect 443604 229018 443786 229254
rect 444022 229018 444204 229254
rect 443604 228934 444204 229018
rect 443604 228698 443786 228934
rect 444022 228698 444204 228934
rect 443604 193254 444204 228698
rect 443604 193018 443786 193254
rect 444022 193018 444204 193254
rect 443604 192934 444204 193018
rect 443604 192698 443786 192934
rect 444022 192698 444204 192934
rect 443604 157254 444204 192698
rect 443604 157018 443786 157254
rect 444022 157018 444204 157254
rect 443604 156934 444204 157018
rect 443604 156698 443786 156934
rect 444022 156698 444204 156934
rect 443604 121254 444204 156698
rect 443604 121018 443786 121254
rect 444022 121018 444204 121254
rect 443604 120934 444204 121018
rect 443604 120698 443786 120934
rect 444022 120698 444204 120934
rect 443604 85254 444204 120698
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7022 425786 -6786
rect 426022 -7022 426204 -6786
rect 425604 -7106 426204 -7022
rect 425604 -7342 425786 -7106
rect 426022 -7342 426204 -7106
rect 425604 -7364 426204 -7342
rect 443604 -5866 444204 12698
rect 450804 705758 451404 705780
rect 450804 705522 450986 705758
rect 451222 705522 451404 705758
rect 450804 705438 451404 705522
rect 450804 705202 450986 705438
rect 451222 705202 451404 705438
rect 450804 668454 451404 705202
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 560454 451404 595898
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 450804 524454 451404 559898
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 450804 488454 451404 523898
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 452454 451404 487898
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 450804 236454 451404 271898
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1266 451404 19898
rect 450804 -1502 450986 -1266
rect 451222 -1502 451404 -1266
rect 450804 -1586 451404 -1502
rect 450804 -1822 450986 -1586
rect 451222 -1822 451404 -1586
rect 450804 -1844 451404 -1822
rect 454404 672054 455004 707042
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 600054 455004 635498
rect 454404 599818 454586 600054
rect 454822 599818 455004 600054
rect 454404 599734 455004 599818
rect 454404 599498 454586 599734
rect 454822 599498 455004 599734
rect 454404 564054 455004 599498
rect 454404 563818 454586 564054
rect 454822 563818 455004 564054
rect 454404 563734 455004 563818
rect 454404 563498 454586 563734
rect 454822 563498 455004 563734
rect 454404 528054 455004 563498
rect 454404 527818 454586 528054
rect 454822 527818 455004 528054
rect 454404 527734 455004 527818
rect 454404 527498 454586 527734
rect 454822 527498 455004 527734
rect 454404 492054 455004 527498
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 456054 455004 491498
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 384054 455004 419498
rect 454404 383818 454586 384054
rect 454822 383818 455004 384054
rect 454404 383734 455004 383818
rect 454404 383498 454586 383734
rect 454822 383498 455004 383734
rect 454404 348054 455004 383498
rect 454404 347818 454586 348054
rect 454822 347818 455004 348054
rect 454404 347734 455004 347818
rect 454404 347498 454586 347734
rect 454822 347498 455004 347734
rect 454404 312054 455004 347498
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 454404 276054 455004 311498
rect 454404 275818 454586 276054
rect 454822 275818 455004 276054
rect 454404 275734 455004 275818
rect 454404 275498 454586 275734
rect 454822 275498 455004 275734
rect 454404 240054 455004 275498
rect 454404 239818 454586 240054
rect 454822 239818 455004 240054
rect 454404 239734 455004 239818
rect 454404 239498 454586 239734
rect 454822 239498 455004 239734
rect 454404 204054 455004 239498
rect 454404 203818 454586 204054
rect 454822 203818 455004 204054
rect 454404 203734 455004 203818
rect 454404 203498 454586 203734
rect 454822 203498 455004 203734
rect 454404 168054 455004 203498
rect 454404 167818 454586 168054
rect 454822 167818 455004 168054
rect 454404 167734 455004 167818
rect 454404 167498 454586 167734
rect 454822 167498 455004 167734
rect 454404 132054 455004 167498
rect 454404 131818 454586 132054
rect 454822 131818 455004 132054
rect 454404 131734 455004 131818
rect 454404 131498 454586 131734
rect 454822 131498 455004 131734
rect 454404 96054 455004 131498
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3106 455004 23498
rect 454404 -3342 454586 -3106
rect 454822 -3342 455004 -3106
rect 454404 -3426 455004 -3342
rect 454404 -3662 454586 -3426
rect 454822 -3662 455004 -3426
rect 454404 -3684 455004 -3662
rect 458004 675654 458604 708882
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 603654 458604 639098
rect 458004 603418 458186 603654
rect 458422 603418 458604 603654
rect 458004 603334 458604 603418
rect 458004 603098 458186 603334
rect 458422 603098 458604 603334
rect 458004 567654 458604 603098
rect 458004 567418 458186 567654
rect 458422 567418 458604 567654
rect 458004 567334 458604 567418
rect 458004 567098 458186 567334
rect 458422 567098 458604 567334
rect 458004 531654 458604 567098
rect 458004 531418 458186 531654
rect 458422 531418 458604 531654
rect 458004 531334 458604 531418
rect 458004 531098 458186 531334
rect 458422 531098 458604 531334
rect 458004 495654 458604 531098
rect 458004 495418 458186 495654
rect 458422 495418 458604 495654
rect 458004 495334 458604 495418
rect 458004 495098 458186 495334
rect 458422 495098 458604 495334
rect 458004 459654 458604 495098
rect 458004 459418 458186 459654
rect 458422 459418 458604 459654
rect 458004 459334 458604 459418
rect 458004 459098 458186 459334
rect 458422 459098 458604 459334
rect 458004 423654 458604 459098
rect 458004 423418 458186 423654
rect 458422 423418 458604 423654
rect 458004 423334 458604 423418
rect 458004 423098 458186 423334
rect 458422 423098 458604 423334
rect 458004 387654 458604 423098
rect 458004 387418 458186 387654
rect 458422 387418 458604 387654
rect 458004 387334 458604 387418
rect 458004 387098 458186 387334
rect 458422 387098 458604 387334
rect 458004 351654 458604 387098
rect 458004 351418 458186 351654
rect 458422 351418 458604 351654
rect 458004 351334 458604 351418
rect 458004 351098 458186 351334
rect 458422 351098 458604 351334
rect 458004 315654 458604 351098
rect 458004 315418 458186 315654
rect 458422 315418 458604 315654
rect 458004 315334 458604 315418
rect 458004 315098 458186 315334
rect 458422 315098 458604 315334
rect 458004 279654 458604 315098
rect 458004 279418 458186 279654
rect 458422 279418 458604 279654
rect 458004 279334 458604 279418
rect 458004 279098 458186 279334
rect 458422 279098 458604 279334
rect 458004 243654 458604 279098
rect 458004 243418 458186 243654
rect 458422 243418 458604 243654
rect 458004 243334 458604 243418
rect 458004 243098 458186 243334
rect 458422 243098 458604 243334
rect 458004 207654 458604 243098
rect 458004 207418 458186 207654
rect 458422 207418 458604 207654
rect 458004 207334 458604 207418
rect 458004 207098 458186 207334
rect 458422 207098 458604 207334
rect 458004 171654 458604 207098
rect 458004 171418 458186 171654
rect 458422 171418 458604 171654
rect 458004 171334 458604 171418
rect 458004 171098 458186 171334
rect 458422 171098 458604 171334
rect 458004 135654 458604 171098
rect 458004 135418 458186 135654
rect 458422 135418 458604 135654
rect 458004 135334 458604 135418
rect 458004 135098 458186 135334
rect 458422 135098 458604 135334
rect 458004 99654 458604 135098
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -4946 458604 27098
rect 458004 -5182 458186 -4946
rect 458422 -5182 458604 -4946
rect 458004 -5266 458604 -5182
rect 458004 -5502 458186 -5266
rect 458422 -5502 458604 -5266
rect 458004 -5524 458604 -5502
rect 461604 679254 462204 710722
rect 479604 710358 480204 711300
rect 479604 710122 479786 710358
rect 480022 710122 480204 710358
rect 479604 710038 480204 710122
rect 479604 709802 479786 710038
rect 480022 709802 480204 710038
rect 476004 708518 476604 709460
rect 476004 708282 476186 708518
rect 476422 708282 476604 708518
rect 476004 708198 476604 708282
rect 476004 707962 476186 708198
rect 476422 707962 476604 708198
rect 472404 706678 473004 707620
rect 472404 706442 472586 706678
rect 472822 706442 473004 706678
rect 472404 706358 473004 706442
rect 472404 706122 472586 706358
rect 472822 706122 473004 706358
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 607254 462204 642698
rect 461604 607018 461786 607254
rect 462022 607018 462204 607254
rect 461604 606934 462204 607018
rect 461604 606698 461786 606934
rect 462022 606698 462204 606934
rect 461604 571254 462204 606698
rect 461604 571018 461786 571254
rect 462022 571018 462204 571254
rect 461604 570934 462204 571018
rect 461604 570698 461786 570934
rect 462022 570698 462204 570934
rect 461604 535254 462204 570698
rect 461604 535018 461786 535254
rect 462022 535018 462204 535254
rect 461604 534934 462204 535018
rect 461604 534698 461786 534934
rect 462022 534698 462204 534934
rect 461604 499254 462204 534698
rect 461604 499018 461786 499254
rect 462022 499018 462204 499254
rect 461604 498934 462204 499018
rect 461604 498698 461786 498934
rect 462022 498698 462204 498934
rect 461604 463254 462204 498698
rect 461604 463018 461786 463254
rect 462022 463018 462204 463254
rect 461604 462934 462204 463018
rect 461604 462698 461786 462934
rect 462022 462698 462204 462934
rect 461604 427254 462204 462698
rect 461604 427018 461786 427254
rect 462022 427018 462204 427254
rect 461604 426934 462204 427018
rect 461604 426698 461786 426934
rect 462022 426698 462204 426934
rect 461604 391254 462204 426698
rect 461604 391018 461786 391254
rect 462022 391018 462204 391254
rect 461604 390934 462204 391018
rect 461604 390698 461786 390934
rect 462022 390698 462204 390934
rect 461604 355254 462204 390698
rect 461604 355018 461786 355254
rect 462022 355018 462204 355254
rect 461604 354934 462204 355018
rect 461604 354698 461786 354934
rect 462022 354698 462204 354934
rect 461604 319254 462204 354698
rect 461604 319018 461786 319254
rect 462022 319018 462204 319254
rect 461604 318934 462204 319018
rect 461604 318698 461786 318934
rect 462022 318698 462204 318934
rect 461604 283254 462204 318698
rect 461604 283018 461786 283254
rect 462022 283018 462204 283254
rect 461604 282934 462204 283018
rect 461604 282698 461786 282934
rect 462022 282698 462204 282934
rect 461604 247254 462204 282698
rect 461604 247018 461786 247254
rect 462022 247018 462204 247254
rect 461604 246934 462204 247018
rect 461604 246698 461786 246934
rect 462022 246698 462204 246934
rect 461604 211254 462204 246698
rect 461604 211018 461786 211254
rect 462022 211018 462204 211254
rect 461604 210934 462204 211018
rect 461604 210698 461786 210934
rect 462022 210698 462204 210934
rect 461604 175254 462204 210698
rect 461604 175018 461786 175254
rect 462022 175018 462204 175254
rect 461604 174934 462204 175018
rect 461604 174698 461786 174934
rect 462022 174698 462204 174934
rect 461604 139254 462204 174698
rect 461604 139018 461786 139254
rect 462022 139018 462204 139254
rect 461604 138934 462204 139018
rect 461604 138698 461786 138934
rect 462022 138698 462204 138934
rect 461604 103254 462204 138698
rect 461604 103018 461786 103254
rect 462022 103018 462204 103254
rect 461604 102934 462204 103018
rect 461604 102698 461786 102934
rect 462022 102698 462204 102934
rect 461604 67254 462204 102698
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6102 443786 -5866
rect 444022 -6102 444204 -5866
rect 443604 -6186 444204 -6102
rect 443604 -6422 443786 -6186
rect 444022 -6422 444204 -6186
rect 443604 -7364 444204 -6422
rect 461604 -6786 462204 30698
rect 468804 704838 469404 705780
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 578454 469404 613898
rect 468804 578218 468986 578454
rect 469222 578218 469404 578454
rect 468804 578134 469404 578218
rect 468804 577898 468986 578134
rect 469222 577898 469404 578134
rect 468804 542454 469404 577898
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1844 469404 -902
rect 472404 690054 473004 706122
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 582054 473004 617498
rect 472404 581818 472586 582054
rect 472822 581818 473004 582054
rect 472404 581734 473004 581818
rect 472404 581498 472586 581734
rect 472822 581498 473004 581734
rect 472404 546054 473004 581498
rect 472404 545818 472586 546054
rect 472822 545818 473004 546054
rect 472404 545734 473004 545818
rect 472404 545498 472586 545734
rect 472822 545498 473004 545734
rect 472404 510054 473004 545498
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 474054 473004 509498
rect 472404 473818 472586 474054
rect 472822 473818 473004 474054
rect 472404 473734 473004 473818
rect 472404 473498 472586 473734
rect 472822 473498 473004 473734
rect 472404 438054 473004 473498
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 402054 473004 437498
rect 472404 401818 472586 402054
rect 472822 401818 473004 402054
rect 472404 401734 473004 401818
rect 472404 401498 472586 401734
rect 472822 401498 473004 401734
rect 472404 366054 473004 401498
rect 472404 365818 472586 366054
rect 472822 365818 473004 366054
rect 472404 365734 473004 365818
rect 472404 365498 472586 365734
rect 472822 365498 473004 365734
rect 472404 330054 473004 365498
rect 472404 329818 472586 330054
rect 472822 329818 473004 330054
rect 472404 329734 473004 329818
rect 472404 329498 472586 329734
rect 472822 329498 473004 329734
rect 472404 294054 473004 329498
rect 472404 293818 472586 294054
rect 472822 293818 473004 294054
rect 472404 293734 473004 293818
rect 472404 293498 472586 293734
rect 472822 293498 473004 293734
rect 472404 258054 473004 293498
rect 472404 257818 472586 258054
rect 472822 257818 473004 258054
rect 472404 257734 473004 257818
rect 472404 257498 472586 257734
rect 472822 257498 473004 257734
rect 472404 222054 473004 257498
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 186054 473004 221498
rect 472404 185818 472586 186054
rect 472822 185818 473004 186054
rect 472404 185734 473004 185818
rect 472404 185498 472586 185734
rect 472822 185498 473004 185734
rect 472404 150054 473004 185498
rect 472404 149818 472586 150054
rect 472822 149818 473004 150054
rect 472404 149734 473004 149818
rect 472404 149498 472586 149734
rect 472822 149498 473004 149734
rect 472404 114054 473004 149498
rect 472404 113818 472586 114054
rect 472822 113818 473004 114054
rect 472404 113734 473004 113818
rect 472404 113498 472586 113734
rect 472822 113498 473004 113734
rect 472404 78054 473004 113498
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2186 473004 5498
rect 472404 -2422 472586 -2186
rect 472822 -2422 473004 -2186
rect 472404 -2506 473004 -2422
rect 472404 -2742 472586 -2506
rect 472822 -2742 473004 -2506
rect 472404 -3684 473004 -2742
rect 476004 693654 476604 707962
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 585654 476604 621098
rect 476004 585418 476186 585654
rect 476422 585418 476604 585654
rect 476004 585334 476604 585418
rect 476004 585098 476186 585334
rect 476422 585098 476604 585334
rect 476004 549654 476604 585098
rect 476004 549418 476186 549654
rect 476422 549418 476604 549654
rect 476004 549334 476604 549418
rect 476004 549098 476186 549334
rect 476422 549098 476604 549334
rect 476004 513654 476604 549098
rect 476004 513418 476186 513654
rect 476422 513418 476604 513654
rect 476004 513334 476604 513418
rect 476004 513098 476186 513334
rect 476422 513098 476604 513334
rect 476004 477654 476604 513098
rect 476004 477418 476186 477654
rect 476422 477418 476604 477654
rect 476004 477334 476604 477418
rect 476004 477098 476186 477334
rect 476422 477098 476604 477334
rect 476004 441654 476604 477098
rect 476004 441418 476186 441654
rect 476422 441418 476604 441654
rect 476004 441334 476604 441418
rect 476004 441098 476186 441334
rect 476422 441098 476604 441334
rect 476004 405654 476604 441098
rect 476004 405418 476186 405654
rect 476422 405418 476604 405654
rect 476004 405334 476604 405418
rect 476004 405098 476186 405334
rect 476422 405098 476604 405334
rect 476004 369654 476604 405098
rect 476004 369418 476186 369654
rect 476422 369418 476604 369654
rect 476004 369334 476604 369418
rect 476004 369098 476186 369334
rect 476422 369098 476604 369334
rect 476004 333654 476604 369098
rect 476004 333418 476186 333654
rect 476422 333418 476604 333654
rect 476004 333334 476604 333418
rect 476004 333098 476186 333334
rect 476422 333098 476604 333334
rect 476004 297654 476604 333098
rect 476004 297418 476186 297654
rect 476422 297418 476604 297654
rect 476004 297334 476604 297418
rect 476004 297098 476186 297334
rect 476422 297098 476604 297334
rect 476004 261654 476604 297098
rect 476004 261418 476186 261654
rect 476422 261418 476604 261654
rect 476004 261334 476604 261418
rect 476004 261098 476186 261334
rect 476422 261098 476604 261334
rect 476004 225654 476604 261098
rect 476004 225418 476186 225654
rect 476422 225418 476604 225654
rect 476004 225334 476604 225418
rect 476004 225098 476186 225334
rect 476422 225098 476604 225334
rect 476004 189654 476604 225098
rect 476004 189418 476186 189654
rect 476422 189418 476604 189654
rect 476004 189334 476604 189418
rect 476004 189098 476186 189334
rect 476422 189098 476604 189334
rect 476004 153654 476604 189098
rect 476004 153418 476186 153654
rect 476422 153418 476604 153654
rect 476004 153334 476604 153418
rect 476004 153098 476186 153334
rect 476422 153098 476604 153334
rect 476004 117654 476604 153098
rect 476004 117418 476186 117654
rect 476422 117418 476604 117654
rect 476004 117334 476604 117418
rect 476004 117098 476186 117334
rect 476422 117098 476604 117334
rect 476004 81654 476604 117098
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4026 476604 9098
rect 476004 -4262 476186 -4026
rect 476422 -4262 476604 -4026
rect 476004 -4346 476604 -4262
rect 476004 -4582 476186 -4346
rect 476422 -4582 476604 -4346
rect 476004 -5524 476604 -4582
rect 479604 697254 480204 709802
rect 497604 711278 498204 711300
rect 497604 711042 497786 711278
rect 498022 711042 498204 711278
rect 497604 710958 498204 711042
rect 497604 710722 497786 710958
rect 498022 710722 498204 710958
rect 494004 709438 494604 709460
rect 494004 709202 494186 709438
rect 494422 709202 494604 709438
rect 494004 709118 494604 709202
rect 494004 708882 494186 709118
rect 494422 708882 494604 709118
rect 490404 707598 491004 707620
rect 490404 707362 490586 707598
rect 490822 707362 491004 707598
rect 490404 707278 491004 707362
rect 490404 707042 490586 707278
rect 490822 707042 491004 707278
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 589254 480204 624698
rect 479604 589018 479786 589254
rect 480022 589018 480204 589254
rect 479604 588934 480204 589018
rect 479604 588698 479786 588934
rect 480022 588698 480204 588934
rect 479604 553254 480204 588698
rect 479604 553018 479786 553254
rect 480022 553018 480204 553254
rect 479604 552934 480204 553018
rect 479604 552698 479786 552934
rect 480022 552698 480204 552934
rect 479604 517254 480204 552698
rect 479604 517018 479786 517254
rect 480022 517018 480204 517254
rect 479604 516934 480204 517018
rect 479604 516698 479786 516934
rect 480022 516698 480204 516934
rect 479604 481254 480204 516698
rect 479604 481018 479786 481254
rect 480022 481018 480204 481254
rect 479604 480934 480204 481018
rect 479604 480698 479786 480934
rect 480022 480698 480204 480934
rect 479604 445254 480204 480698
rect 479604 445018 479786 445254
rect 480022 445018 480204 445254
rect 479604 444934 480204 445018
rect 479604 444698 479786 444934
rect 480022 444698 480204 444934
rect 479604 409254 480204 444698
rect 479604 409018 479786 409254
rect 480022 409018 480204 409254
rect 479604 408934 480204 409018
rect 479604 408698 479786 408934
rect 480022 408698 480204 408934
rect 479604 373254 480204 408698
rect 479604 373018 479786 373254
rect 480022 373018 480204 373254
rect 479604 372934 480204 373018
rect 479604 372698 479786 372934
rect 480022 372698 480204 372934
rect 479604 337254 480204 372698
rect 479604 337018 479786 337254
rect 480022 337018 480204 337254
rect 479604 336934 480204 337018
rect 479604 336698 479786 336934
rect 480022 336698 480204 336934
rect 479604 301254 480204 336698
rect 479604 301018 479786 301254
rect 480022 301018 480204 301254
rect 479604 300934 480204 301018
rect 479604 300698 479786 300934
rect 480022 300698 480204 300934
rect 479604 265254 480204 300698
rect 479604 265018 479786 265254
rect 480022 265018 480204 265254
rect 479604 264934 480204 265018
rect 479604 264698 479786 264934
rect 480022 264698 480204 264934
rect 479604 229254 480204 264698
rect 479604 229018 479786 229254
rect 480022 229018 480204 229254
rect 479604 228934 480204 229018
rect 479604 228698 479786 228934
rect 480022 228698 480204 228934
rect 479604 193254 480204 228698
rect 479604 193018 479786 193254
rect 480022 193018 480204 193254
rect 479604 192934 480204 193018
rect 479604 192698 479786 192934
rect 480022 192698 480204 192934
rect 479604 157254 480204 192698
rect 479604 157018 479786 157254
rect 480022 157018 480204 157254
rect 479604 156934 480204 157018
rect 479604 156698 479786 156934
rect 480022 156698 480204 156934
rect 479604 121254 480204 156698
rect 479604 121018 479786 121254
rect 480022 121018 480204 121254
rect 479604 120934 480204 121018
rect 479604 120698 479786 120934
rect 480022 120698 480204 120934
rect 479604 85254 480204 120698
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 486804 705758 487404 705780
rect 486804 705522 486986 705758
rect 487222 705522 487404 705758
rect 486804 705438 487404 705522
rect 486804 705202 486986 705438
rect 487222 705202 487404 705438
rect 486804 668454 487404 705202
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 560454 487404 595898
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 524454 487404 559898
rect 486804 524218 486986 524454
rect 487222 524218 487404 524454
rect 486804 524134 487404 524218
rect 486804 523898 486986 524134
rect 487222 523898 487404 524134
rect 486804 488454 487404 523898
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 481587 16828 481653 16829
rect 481587 16764 481588 16828
rect 481652 16764 481653 16828
rect 481587 16763 481653 16764
rect 481590 16557 481650 16763
rect 481587 16556 481653 16557
rect 481587 16492 481588 16556
rect 481652 16492 481653 16556
rect 481587 16491 481653 16492
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7022 461786 -6786
rect 462022 -7022 462204 -6786
rect 461604 -7106 462204 -7022
rect 461604 -7342 461786 -7106
rect 462022 -7342 462204 -7106
rect 461604 -7364 462204 -7342
rect 479604 -5866 480204 12698
rect 486804 -1266 487404 19898
rect 486804 -1502 486986 -1266
rect 487222 -1502 487404 -1266
rect 486804 -1586 487404 -1502
rect 486804 -1822 486986 -1586
rect 487222 -1822 487404 -1586
rect 486804 -1844 487404 -1822
rect 490404 672054 491004 707042
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 600054 491004 635498
rect 490404 599818 490586 600054
rect 490822 599818 491004 600054
rect 490404 599734 491004 599818
rect 490404 599498 490586 599734
rect 490822 599498 491004 599734
rect 490404 564054 491004 599498
rect 490404 563818 490586 564054
rect 490822 563818 491004 564054
rect 490404 563734 491004 563818
rect 490404 563498 490586 563734
rect 490822 563498 491004 563734
rect 490404 528054 491004 563498
rect 490404 527818 490586 528054
rect 490822 527818 491004 528054
rect 490404 527734 491004 527818
rect 490404 527498 490586 527734
rect 490822 527498 491004 527734
rect 490404 492054 491004 527498
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 456054 491004 491498
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 384054 491004 419498
rect 490404 383818 490586 384054
rect 490822 383818 491004 384054
rect 490404 383734 491004 383818
rect 490404 383498 490586 383734
rect 490822 383498 491004 383734
rect 490404 348054 491004 383498
rect 490404 347818 490586 348054
rect 490822 347818 491004 348054
rect 490404 347734 491004 347818
rect 490404 347498 490586 347734
rect 490822 347498 491004 347734
rect 490404 312054 491004 347498
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 276054 491004 311498
rect 490404 275818 490586 276054
rect 490822 275818 491004 276054
rect 490404 275734 491004 275818
rect 490404 275498 490586 275734
rect 490822 275498 491004 275734
rect 490404 240054 491004 275498
rect 490404 239818 490586 240054
rect 490822 239818 491004 240054
rect 490404 239734 491004 239818
rect 490404 239498 490586 239734
rect 490822 239498 491004 239734
rect 490404 204054 491004 239498
rect 490404 203818 490586 204054
rect 490822 203818 491004 204054
rect 490404 203734 491004 203818
rect 490404 203498 490586 203734
rect 490822 203498 491004 203734
rect 490404 168054 491004 203498
rect 490404 167818 490586 168054
rect 490822 167818 491004 168054
rect 490404 167734 491004 167818
rect 490404 167498 490586 167734
rect 490822 167498 491004 167734
rect 490404 132054 491004 167498
rect 490404 131818 490586 132054
rect 490822 131818 491004 132054
rect 490404 131734 491004 131818
rect 490404 131498 490586 131734
rect 490822 131498 491004 131734
rect 490404 96054 491004 131498
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3106 491004 23498
rect 490404 -3342 490586 -3106
rect 490822 -3342 491004 -3106
rect 490404 -3426 491004 -3342
rect 490404 -3662 490586 -3426
rect 490822 -3662 491004 -3426
rect 490404 -3684 491004 -3662
rect 494004 675654 494604 708882
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 603654 494604 639098
rect 494004 603418 494186 603654
rect 494422 603418 494604 603654
rect 494004 603334 494604 603418
rect 494004 603098 494186 603334
rect 494422 603098 494604 603334
rect 494004 567654 494604 603098
rect 494004 567418 494186 567654
rect 494422 567418 494604 567654
rect 494004 567334 494604 567418
rect 494004 567098 494186 567334
rect 494422 567098 494604 567334
rect 494004 531654 494604 567098
rect 494004 531418 494186 531654
rect 494422 531418 494604 531654
rect 494004 531334 494604 531418
rect 494004 531098 494186 531334
rect 494422 531098 494604 531334
rect 494004 495654 494604 531098
rect 494004 495418 494186 495654
rect 494422 495418 494604 495654
rect 494004 495334 494604 495418
rect 494004 495098 494186 495334
rect 494422 495098 494604 495334
rect 494004 459654 494604 495098
rect 494004 459418 494186 459654
rect 494422 459418 494604 459654
rect 494004 459334 494604 459418
rect 494004 459098 494186 459334
rect 494422 459098 494604 459334
rect 494004 423654 494604 459098
rect 494004 423418 494186 423654
rect 494422 423418 494604 423654
rect 494004 423334 494604 423418
rect 494004 423098 494186 423334
rect 494422 423098 494604 423334
rect 494004 387654 494604 423098
rect 494004 387418 494186 387654
rect 494422 387418 494604 387654
rect 494004 387334 494604 387418
rect 494004 387098 494186 387334
rect 494422 387098 494604 387334
rect 494004 351654 494604 387098
rect 494004 351418 494186 351654
rect 494422 351418 494604 351654
rect 494004 351334 494604 351418
rect 494004 351098 494186 351334
rect 494422 351098 494604 351334
rect 494004 315654 494604 351098
rect 494004 315418 494186 315654
rect 494422 315418 494604 315654
rect 494004 315334 494604 315418
rect 494004 315098 494186 315334
rect 494422 315098 494604 315334
rect 494004 279654 494604 315098
rect 494004 279418 494186 279654
rect 494422 279418 494604 279654
rect 494004 279334 494604 279418
rect 494004 279098 494186 279334
rect 494422 279098 494604 279334
rect 494004 243654 494604 279098
rect 494004 243418 494186 243654
rect 494422 243418 494604 243654
rect 494004 243334 494604 243418
rect 494004 243098 494186 243334
rect 494422 243098 494604 243334
rect 494004 207654 494604 243098
rect 494004 207418 494186 207654
rect 494422 207418 494604 207654
rect 494004 207334 494604 207418
rect 494004 207098 494186 207334
rect 494422 207098 494604 207334
rect 494004 171654 494604 207098
rect 494004 171418 494186 171654
rect 494422 171418 494604 171654
rect 494004 171334 494604 171418
rect 494004 171098 494186 171334
rect 494422 171098 494604 171334
rect 494004 135654 494604 171098
rect 494004 135418 494186 135654
rect 494422 135418 494604 135654
rect 494004 135334 494604 135418
rect 494004 135098 494186 135334
rect 494422 135098 494604 135334
rect 494004 99654 494604 135098
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -4946 494604 27098
rect 494004 -5182 494186 -4946
rect 494422 -5182 494604 -4946
rect 494004 -5266 494604 -5182
rect 494004 -5502 494186 -5266
rect 494422 -5502 494604 -5266
rect 494004 -5524 494604 -5502
rect 497604 679254 498204 710722
rect 515604 710358 516204 711300
rect 515604 710122 515786 710358
rect 516022 710122 516204 710358
rect 515604 710038 516204 710122
rect 515604 709802 515786 710038
rect 516022 709802 516204 710038
rect 512004 708518 512604 709460
rect 512004 708282 512186 708518
rect 512422 708282 512604 708518
rect 512004 708198 512604 708282
rect 512004 707962 512186 708198
rect 512422 707962 512604 708198
rect 508404 706678 509004 707620
rect 508404 706442 508586 706678
rect 508822 706442 509004 706678
rect 508404 706358 509004 706442
rect 508404 706122 508586 706358
rect 508822 706122 509004 706358
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 607254 498204 642698
rect 497604 607018 497786 607254
rect 498022 607018 498204 607254
rect 497604 606934 498204 607018
rect 497604 606698 497786 606934
rect 498022 606698 498204 606934
rect 497604 571254 498204 606698
rect 497604 571018 497786 571254
rect 498022 571018 498204 571254
rect 497604 570934 498204 571018
rect 497604 570698 497786 570934
rect 498022 570698 498204 570934
rect 497604 535254 498204 570698
rect 497604 535018 497786 535254
rect 498022 535018 498204 535254
rect 497604 534934 498204 535018
rect 497604 534698 497786 534934
rect 498022 534698 498204 534934
rect 497604 499254 498204 534698
rect 497604 499018 497786 499254
rect 498022 499018 498204 499254
rect 497604 498934 498204 499018
rect 497604 498698 497786 498934
rect 498022 498698 498204 498934
rect 497604 463254 498204 498698
rect 497604 463018 497786 463254
rect 498022 463018 498204 463254
rect 497604 462934 498204 463018
rect 497604 462698 497786 462934
rect 498022 462698 498204 462934
rect 497604 427254 498204 462698
rect 497604 427018 497786 427254
rect 498022 427018 498204 427254
rect 497604 426934 498204 427018
rect 497604 426698 497786 426934
rect 498022 426698 498204 426934
rect 497604 391254 498204 426698
rect 497604 391018 497786 391254
rect 498022 391018 498204 391254
rect 497604 390934 498204 391018
rect 497604 390698 497786 390934
rect 498022 390698 498204 390934
rect 497604 355254 498204 390698
rect 497604 355018 497786 355254
rect 498022 355018 498204 355254
rect 497604 354934 498204 355018
rect 497604 354698 497786 354934
rect 498022 354698 498204 354934
rect 497604 319254 498204 354698
rect 497604 319018 497786 319254
rect 498022 319018 498204 319254
rect 497604 318934 498204 319018
rect 497604 318698 497786 318934
rect 498022 318698 498204 318934
rect 497604 283254 498204 318698
rect 497604 283018 497786 283254
rect 498022 283018 498204 283254
rect 497604 282934 498204 283018
rect 497604 282698 497786 282934
rect 498022 282698 498204 282934
rect 497604 247254 498204 282698
rect 497604 247018 497786 247254
rect 498022 247018 498204 247254
rect 497604 246934 498204 247018
rect 497604 246698 497786 246934
rect 498022 246698 498204 246934
rect 497604 211254 498204 246698
rect 497604 211018 497786 211254
rect 498022 211018 498204 211254
rect 497604 210934 498204 211018
rect 497604 210698 497786 210934
rect 498022 210698 498204 210934
rect 497604 175254 498204 210698
rect 497604 175018 497786 175254
rect 498022 175018 498204 175254
rect 497604 174934 498204 175018
rect 497604 174698 497786 174934
rect 498022 174698 498204 174934
rect 497604 139254 498204 174698
rect 497604 139018 497786 139254
rect 498022 139018 498204 139254
rect 497604 138934 498204 139018
rect 497604 138698 497786 138934
rect 498022 138698 498204 138934
rect 497604 103254 498204 138698
rect 497604 103018 497786 103254
rect 498022 103018 498204 103254
rect 497604 102934 498204 103018
rect 497604 102698 497786 102934
rect 498022 102698 498204 102934
rect 497604 67254 498204 102698
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6102 479786 -5866
rect 480022 -6102 480204 -5866
rect 479604 -6186 480204 -6102
rect 479604 -6422 479786 -6186
rect 480022 -6422 480204 -6186
rect 479604 -7364 480204 -6422
rect 497604 -6786 498204 30698
rect 504804 704838 505404 705780
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 502379 17100 502445 17101
rect 502379 17036 502380 17100
rect 502444 17036 502445 17100
rect 502379 17035 502445 17036
rect 502382 16965 502442 17035
rect 502379 16964 502445 16965
rect 502379 16900 502380 16964
rect 502444 16900 502445 16964
rect 502379 16899 502445 16900
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1844 505404 -902
rect 508404 690054 509004 706122
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 546054 509004 581498
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2186 509004 5498
rect 508404 -2422 508586 -2186
rect 508822 -2422 509004 -2186
rect 508404 -2506 509004 -2422
rect 508404 -2742 508586 -2506
rect 508822 -2742 509004 -2506
rect 508404 -3684 509004 -2742
rect 512004 693654 512604 707962
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4026 512604 9098
rect 512004 -4262 512186 -4026
rect 512422 -4262 512604 -4026
rect 512004 -4346 512604 -4262
rect 512004 -4582 512186 -4346
rect 512422 -4582 512604 -4346
rect 512004 -5524 512604 -4582
rect 515604 697254 516204 709802
rect 533604 711278 534204 711300
rect 533604 711042 533786 711278
rect 534022 711042 534204 711278
rect 533604 710958 534204 711042
rect 533604 710722 533786 710958
rect 534022 710722 534204 710958
rect 530004 709438 530604 709460
rect 530004 709202 530186 709438
rect 530422 709202 530604 709438
rect 530004 709118 530604 709202
rect 530004 708882 530186 709118
rect 530422 708882 530604 709118
rect 526404 707598 527004 707620
rect 526404 707362 526586 707598
rect 526822 707362 527004 707598
rect 526404 707278 527004 707362
rect 526404 707042 526586 707278
rect 526822 707042 527004 707278
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7022 497786 -6786
rect 498022 -7022 498204 -6786
rect 497604 -7106 498204 -7022
rect 497604 -7342 497786 -7106
rect 498022 -7342 498204 -7106
rect 497604 -7364 498204 -7342
rect 515604 -5866 516204 12698
rect 522804 705758 523404 705780
rect 522804 705522 522986 705758
rect 523222 705522 523404 705758
rect 522804 705438 523404 705522
rect 522804 705202 522986 705438
rect 523222 705202 523404 705438
rect 522804 668454 523404 705202
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1266 523404 19898
rect 522804 -1502 522986 -1266
rect 523222 -1502 523404 -1266
rect 522804 -1586 523404 -1502
rect 522804 -1822 522986 -1586
rect 523222 -1822 523404 -1586
rect 522804 -1844 523404 -1822
rect 526404 672054 527004 707042
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3106 527004 23498
rect 526404 -3342 526586 -3106
rect 526822 -3342 527004 -3106
rect 526404 -3426 527004 -3342
rect 526404 -3662 526586 -3426
rect 526822 -3662 527004 -3426
rect 526404 -3684 527004 -3662
rect 530004 675654 530604 708882
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -4946 530604 27098
rect 530004 -5182 530186 -4946
rect 530422 -5182 530604 -4946
rect 530004 -5266 530604 -5182
rect 530004 -5502 530186 -5266
rect 530422 -5502 530604 -5266
rect 530004 -5524 530604 -5502
rect 533604 679254 534204 710722
rect 551604 710358 552204 711300
rect 551604 710122 551786 710358
rect 552022 710122 552204 710358
rect 551604 710038 552204 710122
rect 551604 709802 551786 710038
rect 552022 709802 552204 710038
rect 548004 708518 548604 709460
rect 548004 708282 548186 708518
rect 548422 708282 548604 708518
rect 548004 708198 548604 708282
rect 548004 707962 548186 708198
rect 548422 707962 548604 708198
rect 544404 706678 545004 707620
rect 544404 706442 544586 706678
rect 544822 706442 545004 706678
rect 544404 706358 545004 706442
rect 544404 706122 544586 706358
rect 544822 706122 545004 706358
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6102 515786 -5866
rect 516022 -6102 516204 -5866
rect 515604 -6186 516204 -6102
rect 515604 -6422 515786 -6186
rect 516022 -6422 516204 -6186
rect 515604 -7364 516204 -6422
rect 533604 -6786 534204 30698
rect 540804 704838 541404 705780
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1844 541404 -902
rect 544404 690054 545004 706122
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2186 545004 5498
rect 544404 -2422 544586 -2186
rect 544822 -2422 545004 -2186
rect 544404 -2506 545004 -2422
rect 544404 -2742 544586 -2506
rect 544822 -2742 545004 -2506
rect 544404 -3684 545004 -2742
rect 548004 693654 548604 707962
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4026 548604 9098
rect 548004 -4262 548186 -4026
rect 548422 -4262 548604 -4026
rect 548004 -4346 548604 -4262
rect 548004 -4582 548186 -4346
rect 548422 -4582 548604 -4346
rect 548004 -5524 548604 -4582
rect 551604 697254 552204 709802
rect 569604 711278 570204 711300
rect 569604 711042 569786 711278
rect 570022 711042 570204 711278
rect 569604 710958 570204 711042
rect 569604 710722 569786 710958
rect 570022 710722 570204 710958
rect 566004 709438 566604 709460
rect 566004 709202 566186 709438
rect 566422 709202 566604 709438
rect 566004 709118 566604 709202
rect 566004 708882 566186 709118
rect 566422 708882 566604 709118
rect 562404 707598 563004 707620
rect 562404 707362 562586 707598
rect 562822 707362 563004 707598
rect 562404 707278 563004 707362
rect 562404 707042 562586 707278
rect 562822 707042 563004 707278
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7022 533786 -6786
rect 534022 -7022 534204 -6786
rect 533604 -7106 534204 -7022
rect 533604 -7342 533786 -7106
rect 534022 -7342 534204 -7106
rect 533604 -7364 534204 -7342
rect 551604 -5866 552204 12698
rect 558804 705758 559404 705780
rect 558804 705522 558986 705758
rect 559222 705522 559404 705758
rect 558804 705438 559404 705522
rect 558804 705202 558986 705438
rect 559222 705202 559404 705438
rect 558804 668454 559404 705202
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1266 559404 19898
rect 558804 -1502 558986 -1266
rect 559222 -1502 559404 -1266
rect 558804 -1586 559404 -1502
rect 558804 -1822 558986 -1586
rect 559222 -1822 559404 -1586
rect 558804 -1844 559404 -1822
rect 562404 672054 563004 707042
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3106 563004 23498
rect 562404 -3342 562586 -3106
rect 562822 -3342 563004 -3106
rect 562404 -3426 563004 -3342
rect 562404 -3662 562586 -3426
rect 562822 -3662 563004 -3426
rect 562404 -3684 563004 -3662
rect 566004 675654 566604 708882
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -4946 566604 27098
rect 566004 -5182 566186 -4946
rect 566422 -5182 566604 -4946
rect 566004 -5266 566604 -5182
rect 566004 -5502 566186 -5266
rect 566422 -5502 566604 -5266
rect 566004 -5524 566604 -5502
rect 569604 679254 570204 710722
rect 591760 711278 592360 711300
rect 591760 711042 591942 711278
rect 592178 711042 592360 711278
rect 591760 710958 592360 711042
rect 591760 710722 591942 710958
rect 592178 710722 592360 710958
rect 590840 710358 591440 710380
rect 590840 710122 591022 710358
rect 591258 710122 591440 710358
rect 590840 710038 591440 710122
rect 590840 709802 591022 710038
rect 591258 709802 591440 710038
rect 589920 709438 590520 709460
rect 589920 709202 590102 709438
rect 590338 709202 590520 709438
rect 589920 709118 590520 709202
rect 589920 708882 590102 709118
rect 590338 708882 590520 709118
rect 589000 708518 589600 708540
rect 589000 708282 589182 708518
rect 589418 708282 589600 708518
rect 589000 708198 589600 708282
rect 589000 707962 589182 708198
rect 589418 707962 589600 708198
rect 580404 706678 581004 707620
rect 588080 707598 588680 707620
rect 588080 707362 588262 707598
rect 588498 707362 588680 707598
rect 588080 707278 588680 707362
rect 588080 707042 588262 707278
rect 588498 707042 588680 707278
rect 580404 706442 580586 706678
rect 580822 706442 581004 706678
rect 580404 706358 581004 706442
rect 580404 706122 580586 706358
rect 580822 706122 581004 706358
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6102 551786 -5866
rect 552022 -6102 552204 -5866
rect 551604 -6186 552204 -6102
rect 551604 -6422 551786 -6186
rect 552022 -6422 552204 -6186
rect 551604 -7364 552204 -6422
rect 569604 -6786 570204 30698
rect 576804 704838 577404 705780
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1844 577404 -902
rect 580404 690054 581004 706122
rect 587160 706678 587760 706700
rect 587160 706442 587342 706678
rect 587578 706442 587760 706678
rect 587160 706358 587760 706442
rect 587160 706122 587342 706358
rect 587578 706122 587760 706358
rect 586240 705758 586840 705780
rect 586240 705522 586422 705758
rect 586658 705522 586840 705758
rect 586240 705438 586840 705522
rect 586240 705202 586422 705438
rect 586658 705202 586840 705438
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2186 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586240 668454 586840 705202
rect 586240 668218 586422 668454
rect 586658 668218 586840 668454
rect 586240 668134 586840 668218
rect 586240 667898 586422 668134
rect 586658 667898 586840 668134
rect 586240 632454 586840 667898
rect 586240 632218 586422 632454
rect 586658 632218 586840 632454
rect 586240 632134 586840 632218
rect 586240 631898 586422 632134
rect 586658 631898 586840 632134
rect 586240 596454 586840 631898
rect 586240 596218 586422 596454
rect 586658 596218 586840 596454
rect 586240 596134 586840 596218
rect 586240 595898 586422 596134
rect 586658 595898 586840 596134
rect 586240 560454 586840 595898
rect 586240 560218 586422 560454
rect 586658 560218 586840 560454
rect 586240 560134 586840 560218
rect 586240 559898 586422 560134
rect 586658 559898 586840 560134
rect 586240 524454 586840 559898
rect 586240 524218 586422 524454
rect 586658 524218 586840 524454
rect 586240 524134 586840 524218
rect 586240 523898 586422 524134
rect 586658 523898 586840 524134
rect 586240 488454 586840 523898
rect 586240 488218 586422 488454
rect 586658 488218 586840 488454
rect 586240 488134 586840 488218
rect 586240 487898 586422 488134
rect 586658 487898 586840 488134
rect 586240 452454 586840 487898
rect 586240 452218 586422 452454
rect 586658 452218 586840 452454
rect 586240 452134 586840 452218
rect 586240 451898 586422 452134
rect 586658 451898 586840 452134
rect 586240 416454 586840 451898
rect 586240 416218 586422 416454
rect 586658 416218 586840 416454
rect 586240 416134 586840 416218
rect 586240 415898 586422 416134
rect 586658 415898 586840 416134
rect 586240 380454 586840 415898
rect 586240 380218 586422 380454
rect 586658 380218 586840 380454
rect 586240 380134 586840 380218
rect 586240 379898 586422 380134
rect 586658 379898 586840 380134
rect 586240 344454 586840 379898
rect 586240 344218 586422 344454
rect 586658 344218 586840 344454
rect 586240 344134 586840 344218
rect 586240 343898 586422 344134
rect 586658 343898 586840 344134
rect 586240 308454 586840 343898
rect 586240 308218 586422 308454
rect 586658 308218 586840 308454
rect 586240 308134 586840 308218
rect 586240 307898 586422 308134
rect 586658 307898 586840 308134
rect 586240 272454 586840 307898
rect 586240 272218 586422 272454
rect 586658 272218 586840 272454
rect 586240 272134 586840 272218
rect 586240 271898 586422 272134
rect 586658 271898 586840 272134
rect 586240 236454 586840 271898
rect 586240 236218 586422 236454
rect 586658 236218 586840 236454
rect 586240 236134 586840 236218
rect 586240 235898 586422 236134
rect 586658 235898 586840 236134
rect 586240 200454 586840 235898
rect 586240 200218 586422 200454
rect 586658 200218 586840 200454
rect 586240 200134 586840 200218
rect 586240 199898 586422 200134
rect 586658 199898 586840 200134
rect 586240 164454 586840 199898
rect 586240 164218 586422 164454
rect 586658 164218 586840 164454
rect 586240 164134 586840 164218
rect 586240 163898 586422 164134
rect 586658 163898 586840 164134
rect 586240 128454 586840 163898
rect 586240 128218 586422 128454
rect 586658 128218 586840 128454
rect 586240 128134 586840 128218
rect 586240 127898 586422 128134
rect 586658 127898 586840 128134
rect 586240 92454 586840 127898
rect 586240 92218 586422 92454
rect 586658 92218 586840 92454
rect 586240 92134 586840 92218
rect 586240 91898 586422 92134
rect 586658 91898 586840 92134
rect 586240 56454 586840 91898
rect 586240 56218 586422 56454
rect 586658 56218 586840 56454
rect 586240 56134 586840 56218
rect 586240 55898 586422 56134
rect 586658 55898 586840 56134
rect 586240 20454 586840 55898
rect 586240 20218 586422 20454
rect 586658 20218 586840 20454
rect 586240 20134 586840 20218
rect 586240 19898 586422 20134
rect 586658 19898 586840 20134
rect 586240 -1266 586840 19898
rect 586240 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect 586240 -1586 586840 -1502
rect 586240 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect 586240 -1844 586840 -1822
rect 587160 690054 587760 706122
rect 587160 689818 587342 690054
rect 587578 689818 587760 690054
rect 587160 689734 587760 689818
rect 587160 689498 587342 689734
rect 587578 689498 587760 689734
rect 587160 654054 587760 689498
rect 587160 653818 587342 654054
rect 587578 653818 587760 654054
rect 587160 653734 587760 653818
rect 587160 653498 587342 653734
rect 587578 653498 587760 653734
rect 587160 618054 587760 653498
rect 587160 617818 587342 618054
rect 587578 617818 587760 618054
rect 587160 617734 587760 617818
rect 587160 617498 587342 617734
rect 587578 617498 587760 617734
rect 587160 582054 587760 617498
rect 587160 581818 587342 582054
rect 587578 581818 587760 582054
rect 587160 581734 587760 581818
rect 587160 581498 587342 581734
rect 587578 581498 587760 581734
rect 587160 546054 587760 581498
rect 587160 545818 587342 546054
rect 587578 545818 587760 546054
rect 587160 545734 587760 545818
rect 587160 545498 587342 545734
rect 587578 545498 587760 545734
rect 587160 510054 587760 545498
rect 587160 509818 587342 510054
rect 587578 509818 587760 510054
rect 587160 509734 587760 509818
rect 587160 509498 587342 509734
rect 587578 509498 587760 509734
rect 587160 474054 587760 509498
rect 587160 473818 587342 474054
rect 587578 473818 587760 474054
rect 587160 473734 587760 473818
rect 587160 473498 587342 473734
rect 587578 473498 587760 473734
rect 587160 438054 587760 473498
rect 587160 437818 587342 438054
rect 587578 437818 587760 438054
rect 587160 437734 587760 437818
rect 587160 437498 587342 437734
rect 587578 437498 587760 437734
rect 587160 402054 587760 437498
rect 587160 401818 587342 402054
rect 587578 401818 587760 402054
rect 587160 401734 587760 401818
rect 587160 401498 587342 401734
rect 587578 401498 587760 401734
rect 587160 366054 587760 401498
rect 587160 365818 587342 366054
rect 587578 365818 587760 366054
rect 587160 365734 587760 365818
rect 587160 365498 587342 365734
rect 587578 365498 587760 365734
rect 587160 330054 587760 365498
rect 587160 329818 587342 330054
rect 587578 329818 587760 330054
rect 587160 329734 587760 329818
rect 587160 329498 587342 329734
rect 587578 329498 587760 329734
rect 587160 294054 587760 329498
rect 587160 293818 587342 294054
rect 587578 293818 587760 294054
rect 587160 293734 587760 293818
rect 587160 293498 587342 293734
rect 587578 293498 587760 293734
rect 587160 258054 587760 293498
rect 587160 257818 587342 258054
rect 587578 257818 587760 258054
rect 587160 257734 587760 257818
rect 587160 257498 587342 257734
rect 587578 257498 587760 257734
rect 587160 222054 587760 257498
rect 587160 221818 587342 222054
rect 587578 221818 587760 222054
rect 587160 221734 587760 221818
rect 587160 221498 587342 221734
rect 587578 221498 587760 221734
rect 587160 186054 587760 221498
rect 587160 185818 587342 186054
rect 587578 185818 587760 186054
rect 587160 185734 587760 185818
rect 587160 185498 587342 185734
rect 587578 185498 587760 185734
rect 587160 150054 587760 185498
rect 587160 149818 587342 150054
rect 587578 149818 587760 150054
rect 587160 149734 587760 149818
rect 587160 149498 587342 149734
rect 587578 149498 587760 149734
rect 587160 114054 587760 149498
rect 587160 113818 587342 114054
rect 587578 113818 587760 114054
rect 587160 113734 587760 113818
rect 587160 113498 587342 113734
rect 587578 113498 587760 113734
rect 587160 78054 587760 113498
rect 587160 77818 587342 78054
rect 587578 77818 587760 78054
rect 587160 77734 587760 77818
rect 587160 77498 587342 77734
rect 587578 77498 587760 77734
rect 587160 42054 587760 77498
rect 587160 41818 587342 42054
rect 587578 41818 587760 42054
rect 587160 41734 587760 41818
rect 587160 41498 587342 41734
rect 587578 41498 587760 41734
rect 587160 6054 587760 41498
rect 587160 5818 587342 6054
rect 587578 5818 587760 6054
rect 587160 5734 587760 5818
rect 587160 5498 587342 5734
rect 587578 5498 587760 5734
rect 580404 -2422 580586 -2186
rect 580822 -2422 581004 -2186
rect 580404 -2506 581004 -2422
rect 580404 -2742 580586 -2506
rect 580822 -2742 581004 -2506
rect 580404 -3684 581004 -2742
rect 587160 -2186 587760 5498
rect 587160 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect 587160 -2506 587760 -2422
rect 587160 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect 587160 -2764 587760 -2742
rect 588080 672054 588680 707042
rect 588080 671818 588262 672054
rect 588498 671818 588680 672054
rect 588080 671734 588680 671818
rect 588080 671498 588262 671734
rect 588498 671498 588680 671734
rect 588080 636054 588680 671498
rect 588080 635818 588262 636054
rect 588498 635818 588680 636054
rect 588080 635734 588680 635818
rect 588080 635498 588262 635734
rect 588498 635498 588680 635734
rect 588080 600054 588680 635498
rect 588080 599818 588262 600054
rect 588498 599818 588680 600054
rect 588080 599734 588680 599818
rect 588080 599498 588262 599734
rect 588498 599498 588680 599734
rect 588080 564054 588680 599498
rect 588080 563818 588262 564054
rect 588498 563818 588680 564054
rect 588080 563734 588680 563818
rect 588080 563498 588262 563734
rect 588498 563498 588680 563734
rect 588080 528054 588680 563498
rect 588080 527818 588262 528054
rect 588498 527818 588680 528054
rect 588080 527734 588680 527818
rect 588080 527498 588262 527734
rect 588498 527498 588680 527734
rect 588080 492054 588680 527498
rect 588080 491818 588262 492054
rect 588498 491818 588680 492054
rect 588080 491734 588680 491818
rect 588080 491498 588262 491734
rect 588498 491498 588680 491734
rect 588080 456054 588680 491498
rect 588080 455818 588262 456054
rect 588498 455818 588680 456054
rect 588080 455734 588680 455818
rect 588080 455498 588262 455734
rect 588498 455498 588680 455734
rect 588080 420054 588680 455498
rect 588080 419818 588262 420054
rect 588498 419818 588680 420054
rect 588080 419734 588680 419818
rect 588080 419498 588262 419734
rect 588498 419498 588680 419734
rect 588080 384054 588680 419498
rect 588080 383818 588262 384054
rect 588498 383818 588680 384054
rect 588080 383734 588680 383818
rect 588080 383498 588262 383734
rect 588498 383498 588680 383734
rect 588080 348054 588680 383498
rect 588080 347818 588262 348054
rect 588498 347818 588680 348054
rect 588080 347734 588680 347818
rect 588080 347498 588262 347734
rect 588498 347498 588680 347734
rect 588080 312054 588680 347498
rect 588080 311818 588262 312054
rect 588498 311818 588680 312054
rect 588080 311734 588680 311818
rect 588080 311498 588262 311734
rect 588498 311498 588680 311734
rect 588080 276054 588680 311498
rect 588080 275818 588262 276054
rect 588498 275818 588680 276054
rect 588080 275734 588680 275818
rect 588080 275498 588262 275734
rect 588498 275498 588680 275734
rect 588080 240054 588680 275498
rect 588080 239818 588262 240054
rect 588498 239818 588680 240054
rect 588080 239734 588680 239818
rect 588080 239498 588262 239734
rect 588498 239498 588680 239734
rect 588080 204054 588680 239498
rect 588080 203818 588262 204054
rect 588498 203818 588680 204054
rect 588080 203734 588680 203818
rect 588080 203498 588262 203734
rect 588498 203498 588680 203734
rect 588080 168054 588680 203498
rect 588080 167818 588262 168054
rect 588498 167818 588680 168054
rect 588080 167734 588680 167818
rect 588080 167498 588262 167734
rect 588498 167498 588680 167734
rect 588080 132054 588680 167498
rect 588080 131818 588262 132054
rect 588498 131818 588680 132054
rect 588080 131734 588680 131818
rect 588080 131498 588262 131734
rect 588498 131498 588680 131734
rect 588080 96054 588680 131498
rect 588080 95818 588262 96054
rect 588498 95818 588680 96054
rect 588080 95734 588680 95818
rect 588080 95498 588262 95734
rect 588498 95498 588680 95734
rect 588080 60054 588680 95498
rect 588080 59818 588262 60054
rect 588498 59818 588680 60054
rect 588080 59734 588680 59818
rect 588080 59498 588262 59734
rect 588498 59498 588680 59734
rect 588080 24054 588680 59498
rect 588080 23818 588262 24054
rect 588498 23818 588680 24054
rect 588080 23734 588680 23818
rect 588080 23498 588262 23734
rect 588498 23498 588680 23734
rect 588080 -3106 588680 23498
rect 588080 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect 588080 -3426 588680 -3342
rect 588080 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect 588080 -3684 588680 -3662
rect 589000 693654 589600 707962
rect 589000 693418 589182 693654
rect 589418 693418 589600 693654
rect 589000 693334 589600 693418
rect 589000 693098 589182 693334
rect 589418 693098 589600 693334
rect 589000 657654 589600 693098
rect 589000 657418 589182 657654
rect 589418 657418 589600 657654
rect 589000 657334 589600 657418
rect 589000 657098 589182 657334
rect 589418 657098 589600 657334
rect 589000 621654 589600 657098
rect 589000 621418 589182 621654
rect 589418 621418 589600 621654
rect 589000 621334 589600 621418
rect 589000 621098 589182 621334
rect 589418 621098 589600 621334
rect 589000 585654 589600 621098
rect 589000 585418 589182 585654
rect 589418 585418 589600 585654
rect 589000 585334 589600 585418
rect 589000 585098 589182 585334
rect 589418 585098 589600 585334
rect 589000 549654 589600 585098
rect 589000 549418 589182 549654
rect 589418 549418 589600 549654
rect 589000 549334 589600 549418
rect 589000 549098 589182 549334
rect 589418 549098 589600 549334
rect 589000 513654 589600 549098
rect 589000 513418 589182 513654
rect 589418 513418 589600 513654
rect 589000 513334 589600 513418
rect 589000 513098 589182 513334
rect 589418 513098 589600 513334
rect 589000 477654 589600 513098
rect 589000 477418 589182 477654
rect 589418 477418 589600 477654
rect 589000 477334 589600 477418
rect 589000 477098 589182 477334
rect 589418 477098 589600 477334
rect 589000 441654 589600 477098
rect 589000 441418 589182 441654
rect 589418 441418 589600 441654
rect 589000 441334 589600 441418
rect 589000 441098 589182 441334
rect 589418 441098 589600 441334
rect 589000 405654 589600 441098
rect 589000 405418 589182 405654
rect 589418 405418 589600 405654
rect 589000 405334 589600 405418
rect 589000 405098 589182 405334
rect 589418 405098 589600 405334
rect 589000 369654 589600 405098
rect 589000 369418 589182 369654
rect 589418 369418 589600 369654
rect 589000 369334 589600 369418
rect 589000 369098 589182 369334
rect 589418 369098 589600 369334
rect 589000 333654 589600 369098
rect 589000 333418 589182 333654
rect 589418 333418 589600 333654
rect 589000 333334 589600 333418
rect 589000 333098 589182 333334
rect 589418 333098 589600 333334
rect 589000 297654 589600 333098
rect 589000 297418 589182 297654
rect 589418 297418 589600 297654
rect 589000 297334 589600 297418
rect 589000 297098 589182 297334
rect 589418 297098 589600 297334
rect 589000 261654 589600 297098
rect 589000 261418 589182 261654
rect 589418 261418 589600 261654
rect 589000 261334 589600 261418
rect 589000 261098 589182 261334
rect 589418 261098 589600 261334
rect 589000 225654 589600 261098
rect 589000 225418 589182 225654
rect 589418 225418 589600 225654
rect 589000 225334 589600 225418
rect 589000 225098 589182 225334
rect 589418 225098 589600 225334
rect 589000 189654 589600 225098
rect 589000 189418 589182 189654
rect 589418 189418 589600 189654
rect 589000 189334 589600 189418
rect 589000 189098 589182 189334
rect 589418 189098 589600 189334
rect 589000 153654 589600 189098
rect 589000 153418 589182 153654
rect 589418 153418 589600 153654
rect 589000 153334 589600 153418
rect 589000 153098 589182 153334
rect 589418 153098 589600 153334
rect 589000 117654 589600 153098
rect 589000 117418 589182 117654
rect 589418 117418 589600 117654
rect 589000 117334 589600 117418
rect 589000 117098 589182 117334
rect 589418 117098 589600 117334
rect 589000 81654 589600 117098
rect 589000 81418 589182 81654
rect 589418 81418 589600 81654
rect 589000 81334 589600 81418
rect 589000 81098 589182 81334
rect 589418 81098 589600 81334
rect 589000 45654 589600 81098
rect 589000 45418 589182 45654
rect 589418 45418 589600 45654
rect 589000 45334 589600 45418
rect 589000 45098 589182 45334
rect 589418 45098 589600 45334
rect 589000 9654 589600 45098
rect 589000 9418 589182 9654
rect 589418 9418 589600 9654
rect 589000 9334 589600 9418
rect 589000 9098 589182 9334
rect 589418 9098 589600 9334
rect 589000 -4026 589600 9098
rect 589000 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect 589000 -4346 589600 -4262
rect 589000 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect 589000 -4604 589600 -4582
rect 589920 675654 590520 708882
rect 589920 675418 590102 675654
rect 590338 675418 590520 675654
rect 589920 675334 590520 675418
rect 589920 675098 590102 675334
rect 590338 675098 590520 675334
rect 589920 639654 590520 675098
rect 589920 639418 590102 639654
rect 590338 639418 590520 639654
rect 589920 639334 590520 639418
rect 589920 639098 590102 639334
rect 590338 639098 590520 639334
rect 589920 603654 590520 639098
rect 589920 603418 590102 603654
rect 590338 603418 590520 603654
rect 589920 603334 590520 603418
rect 589920 603098 590102 603334
rect 590338 603098 590520 603334
rect 589920 567654 590520 603098
rect 589920 567418 590102 567654
rect 590338 567418 590520 567654
rect 589920 567334 590520 567418
rect 589920 567098 590102 567334
rect 590338 567098 590520 567334
rect 589920 531654 590520 567098
rect 589920 531418 590102 531654
rect 590338 531418 590520 531654
rect 589920 531334 590520 531418
rect 589920 531098 590102 531334
rect 590338 531098 590520 531334
rect 589920 495654 590520 531098
rect 589920 495418 590102 495654
rect 590338 495418 590520 495654
rect 589920 495334 590520 495418
rect 589920 495098 590102 495334
rect 590338 495098 590520 495334
rect 589920 459654 590520 495098
rect 589920 459418 590102 459654
rect 590338 459418 590520 459654
rect 589920 459334 590520 459418
rect 589920 459098 590102 459334
rect 590338 459098 590520 459334
rect 589920 423654 590520 459098
rect 589920 423418 590102 423654
rect 590338 423418 590520 423654
rect 589920 423334 590520 423418
rect 589920 423098 590102 423334
rect 590338 423098 590520 423334
rect 589920 387654 590520 423098
rect 589920 387418 590102 387654
rect 590338 387418 590520 387654
rect 589920 387334 590520 387418
rect 589920 387098 590102 387334
rect 590338 387098 590520 387334
rect 589920 351654 590520 387098
rect 589920 351418 590102 351654
rect 590338 351418 590520 351654
rect 589920 351334 590520 351418
rect 589920 351098 590102 351334
rect 590338 351098 590520 351334
rect 589920 315654 590520 351098
rect 589920 315418 590102 315654
rect 590338 315418 590520 315654
rect 589920 315334 590520 315418
rect 589920 315098 590102 315334
rect 590338 315098 590520 315334
rect 589920 279654 590520 315098
rect 589920 279418 590102 279654
rect 590338 279418 590520 279654
rect 589920 279334 590520 279418
rect 589920 279098 590102 279334
rect 590338 279098 590520 279334
rect 589920 243654 590520 279098
rect 589920 243418 590102 243654
rect 590338 243418 590520 243654
rect 589920 243334 590520 243418
rect 589920 243098 590102 243334
rect 590338 243098 590520 243334
rect 589920 207654 590520 243098
rect 589920 207418 590102 207654
rect 590338 207418 590520 207654
rect 589920 207334 590520 207418
rect 589920 207098 590102 207334
rect 590338 207098 590520 207334
rect 589920 171654 590520 207098
rect 589920 171418 590102 171654
rect 590338 171418 590520 171654
rect 589920 171334 590520 171418
rect 589920 171098 590102 171334
rect 590338 171098 590520 171334
rect 589920 135654 590520 171098
rect 589920 135418 590102 135654
rect 590338 135418 590520 135654
rect 589920 135334 590520 135418
rect 589920 135098 590102 135334
rect 590338 135098 590520 135334
rect 589920 99654 590520 135098
rect 589920 99418 590102 99654
rect 590338 99418 590520 99654
rect 589920 99334 590520 99418
rect 589920 99098 590102 99334
rect 590338 99098 590520 99334
rect 589920 63654 590520 99098
rect 589920 63418 590102 63654
rect 590338 63418 590520 63654
rect 589920 63334 590520 63418
rect 589920 63098 590102 63334
rect 590338 63098 590520 63334
rect 589920 27654 590520 63098
rect 589920 27418 590102 27654
rect 590338 27418 590520 27654
rect 589920 27334 590520 27418
rect 589920 27098 590102 27334
rect 590338 27098 590520 27334
rect 589920 -4946 590520 27098
rect 589920 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect 589920 -5266 590520 -5182
rect 589920 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect 589920 -5524 590520 -5502
rect 590840 697254 591440 709802
rect 590840 697018 591022 697254
rect 591258 697018 591440 697254
rect 590840 696934 591440 697018
rect 590840 696698 591022 696934
rect 591258 696698 591440 696934
rect 590840 661254 591440 696698
rect 590840 661018 591022 661254
rect 591258 661018 591440 661254
rect 590840 660934 591440 661018
rect 590840 660698 591022 660934
rect 591258 660698 591440 660934
rect 590840 625254 591440 660698
rect 590840 625018 591022 625254
rect 591258 625018 591440 625254
rect 590840 624934 591440 625018
rect 590840 624698 591022 624934
rect 591258 624698 591440 624934
rect 590840 589254 591440 624698
rect 590840 589018 591022 589254
rect 591258 589018 591440 589254
rect 590840 588934 591440 589018
rect 590840 588698 591022 588934
rect 591258 588698 591440 588934
rect 590840 553254 591440 588698
rect 590840 553018 591022 553254
rect 591258 553018 591440 553254
rect 590840 552934 591440 553018
rect 590840 552698 591022 552934
rect 591258 552698 591440 552934
rect 590840 517254 591440 552698
rect 590840 517018 591022 517254
rect 591258 517018 591440 517254
rect 590840 516934 591440 517018
rect 590840 516698 591022 516934
rect 591258 516698 591440 516934
rect 590840 481254 591440 516698
rect 590840 481018 591022 481254
rect 591258 481018 591440 481254
rect 590840 480934 591440 481018
rect 590840 480698 591022 480934
rect 591258 480698 591440 480934
rect 590840 445254 591440 480698
rect 590840 445018 591022 445254
rect 591258 445018 591440 445254
rect 590840 444934 591440 445018
rect 590840 444698 591022 444934
rect 591258 444698 591440 444934
rect 590840 409254 591440 444698
rect 590840 409018 591022 409254
rect 591258 409018 591440 409254
rect 590840 408934 591440 409018
rect 590840 408698 591022 408934
rect 591258 408698 591440 408934
rect 590840 373254 591440 408698
rect 590840 373018 591022 373254
rect 591258 373018 591440 373254
rect 590840 372934 591440 373018
rect 590840 372698 591022 372934
rect 591258 372698 591440 372934
rect 590840 337254 591440 372698
rect 590840 337018 591022 337254
rect 591258 337018 591440 337254
rect 590840 336934 591440 337018
rect 590840 336698 591022 336934
rect 591258 336698 591440 336934
rect 590840 301254 591440 336698
rect 590840 301018 591022 301254
rect 591258 301018 591440 301254
rect 590840 300934 591440 301018
rect 590840 300698 591022 300934
rect 591258 300698 591440 300934
rect 590840 265254 591440 300698
rect 590840 265018 591022 265254
rect 591258 265018 591440 265254
rect 590840 264934 591440 265018
rect 590840 264698 591022 264934
rect 591258 264698 591440 264934
rect 590840 229254 591440 264698
rect 590840 229018 591022 229254
rect 591258 229018 591440 229254
rect 590840 228934 591440 229018
rect 590840 228698 591022 228934
rect 591258 228698 591440 228934
rect 590840 193254 591440 228698
rect 590840 193018 591022 193254
rect 591258 193018 591440 193254
rect 590840 192934 591440 193018
rect 590840 192698 591022 192934
rect 591258 192698 591440 192934
rect 590840 157254 591440 192698
rect 590840 157018 591022 157254
rect 591258 157018 591440 157254
rect 590840 156934 591440 157018
rect 590840 156698 591022 156934
rect 591258 156698 591440 156934
rect 590840 121254 591440 156698
rect 590840 121018 591022 121254
rect 591258 121018 591440 121254
rect 590840 120934 591440 121018
rect 590840 120698 591022 120934
rect 591258 120698 591440 120934
rect 590840 85254 591440 120698
rect 590840 85018 591022 85254
rect 591258 85018 591440 85254
rect 590840 84934 591440 85018
rect 590840 84698 591022 84934
rect 591258 84698 591440 84934
rect 590840 49254 591440 84698
rect 590840 49018 591022 49254
rect 591258 49018 591440 49254
rect 590840 48934 591440 49018
rect 590840 48698 591022 48934
rect 591258 48698 591440 48934
rect 590840 13254 591440 48698
rect 590840 13018 591022 13254
rect 591258 13018 591440 13254
rect 590840 12934 591440 13018
rect 590840 12698 591022 12934
rect 591258 12698 591440 12934
rect 590840 -5866 591440 12698
rect 590840 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect 590840 -6186 591440 -6102
rect 590840 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect 590840 -6444 591440 -6422
rect 591760 679254 592360 710722
rect 591760 679018 591942 679254
rect 592178 679018 592360 679254
rect 591760 678934 592360 679018
rect 591760 678698 591942 678934
rect 592178 678698 592360 678934
rect 591760 643254 592360 678698
rect 591760 643018 591942 643254
rect 592178 643018 592360 643254
rect 591760 642934 592360 643018
rect 591760 642698 591942 642934
rect 592178 642698 592360 642934
rect 591760 607254 592360 642698
rect 591760 607018 591942 607254
rect 592178 607018 592360 607254
rect 591760 606934 592360 607018
rect 591760 606698 591942 606934
rect 592178 606698 592360 606934
rect 591760 571254 592360 606698
rect 591760 571018 591942 571254
rect 592178 571018 592360 571254
rect 591760 570934 592360 571018
rect 591760 570698 591942 570934
rect 592178 570698 592360 570934
rect 591760 535254 592360 570698
rect 591760 535018 591942 535254
rect 592178 535018 592360 535254
rect 591760 534934 592360 535018
rect 591760 534698 591942 534934
rect 592178 534698 592360 534934
rect 591760 499254 592360 534698
rect 591760 499018 591942 499254
rect 592178 499018 592360 499254
rect 591760 498934 592360 499018
rect 591760 498698 591942 498934
rect 592178 498698 592360 498934
rect 591760 463254 592360 498698
rect 591760 463018 591942 463254
rect 592178 463018 592360 463254
rect 591760 462934 592360 463018
rect 591760 462698 591942 462934
rect 592178 462698 592360 462934
rect 591760 427254 592360 462698
rect 591760 427018 591942 427254
rect 592178 427018 592360 427254
rect 591760 426934 592360 427018
rect 591760 426698 591942 426934
rect 592178 426698 592360 426934
rect 591760 391254 592360 426698
rect 591760 391018 591942 391254
rect 592178 391018 592360 391254
rect 591760 390934 592360 391018
rect 591760 390698 591942 390934
rect 592178 390698 592360 390934
rect 591760 355254 592360 390698
rect 591760 355018 591942 355254
rect 592178 355018 592360 355254
rect 591760 354934 592360 355018
rect 591760 354698 591942 354934
rect 592178 354698 592360 354934
rect 591760 319254 592360 354698
rect 591760 319018 591942 319254
rect 592178 319018 592360 319254
rect 591760 318934 592360 319018
rect 591760 318698 591942 318934
rect 592178 318698 592360 318934
rect 591760 283254 592360 318698
rect 591760 283018 591942 283254
rect 592178 283018 592360 283254
rect 591760 282934 592360 283018
rect 591760 282698 591942 282934
rect 592178 282698 592360 282934
rect 591760 247254 592360 282698
rect 591760 247018 591942 247254
rect 592178 247018 592360 247254
rect 591760 246934 592360 247018
rect 591760 246698 591942 246934
rect 592178 246698 592360 246934
rect 591760 211254 592360 246698
rect 591760 211018 591942 211254
rect 592178 211018 592360 211254
rect 591760 210934 592360 211018
rect 591760 210698 591942 210934
rect 592178 210698 592360 210934
rect 591760 175254 592360 210698
rect 591760 175018 591942 175254
rect 592178 175018 592360 175254
rect 591760 174934 592360 175018
rect 591760 174698 591942 174934
rect 592178 174698 592360 174934
rect 591760 139254 592360 174698
rect 591760 139018 591942 139254
rect 592178 139018 592360 139254
rect 591760 138934 592360 139018
rect 591760 138698 591942 138934
rect 592178 138698 592360 138934
rect 591760 103254 592360 138698
rect 591760 103018 591942 103254
rect 592178 103018 592360 103254
rect 591760 102934 592360 103018
rect 591760 102698 591942 102934
rect 592178 102698 592360 102934
rect 591760 67254 592360 102698
rect 591760 67018 591942 67254
rect 592178 67018 592360 67254
rect 591760 66934 592360 67018
rect 591760 66698 591942 66934
rect 592178 66698 592360 66934
rect 591760 31254 592360 66698
rect 591760 31018 591942 31254
rect 592178 31018 592360 31254
rect 591760 30934 592360 31018
rect 591760 30698 591942 30934
rect 592178 30698 592360 30934
rect 569604 -7022 569786 -6786
rect 570022 -7022 570204 -6786
rect 569604 -7106 570204 -7022
rect 569604 -7342 569786 -7106
rect 570022 -7342 570204 -7106
rect 569604 -7364 570204 -7342
rect 591760 -6786 592360 30698
rect 591760 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect 591760 -7106 592360 -7022
rect 591760 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect 591760 -7364 592360 -7342
<< via4 >>
rect -8254 711042 -8018 711278
rect -8254 710722 -8018 710958
rect -8254 679018 -8018 679254
rect -8254 678698 -8018 678934
rect -8254 643018 -8018 643254
rect -8254 642698 -8018 642934
rect -8254 607018 -8018 607254
rect -8254 606698 -8018 606934
rect -8254 571018 -8018 571254
rect -8254 570698 -8018 570934
rect -8254 535018 -8018 535254
rect -8254 534698 -8018 534934
rect -8254 499018 -8018 499254
rect -8254 498698 -8018 498934
rect -8254 463018 -8018 463254
rect -8254 462698 -8018 462934
rect -8254 427018 -8018 427254
rect -8254 426698 -8018 426934
rect -8254 391018 -8018 391254
rect -8254 390698 -8018 390934
rect -8254 355018 -8018 355254
rect -8254 354698 -8018 354934
rect -8254 319018 -8018 319254
rect -8254 318698 -8018 318934
rect -8254 283018 -8018 283254
rect -8254 282698 -8018 282934
rect -8254 247018 -8018 247254
rect -8254 246698 -8018 246934
rect -8254 211018 -8018 211254
rect -8254 210698 -8018 210934
rect -8254 175018 -8018 175254
rect -8254 174698 -8018 174934
rect -8254 139018 -8018 139254
rect -8254 138698 -8018 138934
rect -8254 103018 -8018 103254
rect -8254 102698 -8018 102934
rect -8254 67018 -8018 67254
rect -8254 66698 -8018 66934
rect -8254 31018 -8018 31254
rect -8254 30698 -8018 30934
rect -7334 710122 -7098 710358
rect -7334 709802 -7098 710038
rect 11786 710122 12022 710358
rect 11786 709802 12022 710038
rect -7334 697018 -7098 697254
rect -7334 696698 -7098 696934
rect -7334 661018 -7098 661254
rect -7334 660698 -7098 660934
rect -7334 625018 -7098 625254
rect -7334 624698 -7098 624934
rect -7334 589018 -7098 589254
rect -7334 588698 -7098 588934
rect -7334 553018 -7098 553254
rect -7334 552698 -7098 552934
rect -7334 517018 -7098 517254
rect -7334 516698 -7098 516934
rect -7334 481018 -7098 481254
rect -7334 480698 -7098 480934
rect -7334 445018 -7098 445254
rect -7334 444698 -7098 444934
rect -7334 409018 -7098 409254
rect -7334 408698 -7098 408934
rect -7334 373018 -7098 373254
rect -7334 372698 -7098 372934
rect -7334 337018 -7098 337254
rect -7334 336698 -7098 336934
rect -7334 301018 -7098 301254
rect -7334 300698 -7098 300934
rect -7334 265018 -7098 265254
rect -7334 264698 -7098 264934
rect -7334 229018 -7098 229254
rect -7334 228698 -7098 228934
rect -7334 193018 -7098 193254
rect -7334 192698 -7098 192934
rect -7334 157018 -7098 157254
rect -7334 156698 -7098 156934
rect -7334 121018 -7098 121254
rect -7334 120698 -7098 120934
rect -7334 85018 -7098 85254
rect -7334 84698 -7098 84934
rect -7334 49018 -7098 49254
rect -7334 48698 -7098 48934
rect -7334 13018 -7098 13254
rect -7334 12698 -7098 12934
rect -6414 709202 -6178 709438
rect -6414 708882 -6178 709118
rect -6414 675418 -6178 675654
rect -6414 675098 -6178 675334
rect -6414 639418 -6178 639654
rect -6414 639098 -6178 639334
rect -6414 603418 -6178 603654
rect -6414 603098 -6178 603334
rect -6414 567418 -6178 567654
rect -6414 567098 -6178 567334
rect -6414 531418 -6178 531654
rect -6414 531098 -6178 531334
rect -6414 495418 -6178 495654
rect -6414 495098 -6178 495334
rect -6414 459418 -6178 459654
rect -6414 459098 -6178 459334
rect -6414 423418 -6178 423654
rect -6414 423098 -6178 423334
rect -6414 387418 -6178 387654
rect -6414 387098 -6178 387334
rect -6414 351418 -6178 351654
rect -6414 351098 -6178 351334
rect -6414 315418 -6178 315654
rect -6414 315098 -6178 315334
rect -6414 279418 -6178 279654
rect -6414 279098 -6178 279334
rect -6414 243418 -6178 243654
rect -6414 243098 -6178 243334
rect -6414 207418 -6178 207654
rect -6414 207098 -6178 207334
rect -6414 171418 -6178 171654
rect -6414 171098 -6178 171334
rect -6414 135418 -6178 135654
rect -6414 135098 -6178 135334
rect -6414 99418 -6178 99654
rect -6414 99098 -6178 99334
rect -6414 63418 -6178 63654
rect -6414 63098 -6178 63334
rect -6414 27418 -6178 27654
rect -6414 27098 -6178 27334
rect -5494 708282 -5258 708518
rect -5494 707962 -5258 708198
rect 8186 708282 8422 708518
rect 8186 707962 8422 708198
rect -5494 693418 -5258 693654
rect -5494 693098 -5258 693334
rect -5494 657418 -5258 657654
rect -5494 657098 -5258 657334
rect -5494 621418 -5258 621654
rect -5494 621098 -5258 621334
rect -5494 585418 -5258 585654
rect -5494 585098 -5258 585334
rect -5494 549418 -5258 549654
rect -5494 549098 -5258 549334
rect -5494 513418 -5258 513654
rect -5494 513098 -5258 513334
rect -5494 477418 -5258 477654
rect -5494 477098 -5258 477334
rect -5494 441418 -5258 441654
rect -5494 441098 -5258 441334
rect -5494 405418 -5258 405654
rect -5494 405098 -5258 405334
rect -5494 369418 -5258 369654
rect -5494 369098 -5258 369334
rect -5494 333418 -5258 333654
rect -5494 333098 -5258 333334
rect -5494 297418 -5258 297654
rect -5494 297098 -5258 297334
rect -5494 261418 -5258 261654
rect -5494 261098 -5258 261334
rect -5494 225418 -5258 225654
rect -5494 225098 -5258 225334
rect -5494 189418 -5258 189654
rect -5494 189098 -5258 189334
rect -5494 153418 -5258 153654
rect -5494 153098 -5258 153334
rect -5494 117418 -5258 117654
rect -5494 117098 -5258 117334
rect -5494 81418 -5258 81654
rect -5494 81098 -5258 81334
rect -5494 45418 -5258 45654
rect -5494 45098 -5258 45334
rect -5494 9418 -5258 9654
rect -5494 9098 -5258 9334
rect -4574 707362 -4338 707598
rect -4574 707042 -4338 707278
rect -4574 671818 -4338 672054
rect -4574 671498 -4338 671734
rect -4574 635818 -4338 636054
rect -4574 635498 -4338 635734
rect -4574 599818 -4338 600054
rect -4574 599498 -4338 599734
rect -4574 563818 -4338 564054
rect -4574 563498 -4338 563734
rect -4574 527818 -4338 528054
rect -4574 527498 -4338 527734
rect -4574 491818 -4338 492054
rect -4574 491498 -4338 491734
rect -4574 455818 -4338 456054
rect -4574 455498 -4338 455734
rect -4574 419818 -4338 420054
rect -4574 419498 -4338 419734
rect -4574 383818 -4338 384054
rect -4574 383498 -4338 383734
rect -4574 347818 -4338 348054
rect -4574 347498 -4338 347734
rect -4574 311818 -4338 312054
rect -4574 311498 -4338 311734
rect -4574 275818 -4338 276054
rect -4574 275498 -4338 275734
rect -4574 239818 -4338 240054
rect -4574 239498 -4338 239734
rect -4574 203818 -4338 204054
rect -4574 203498 -4338 203734
rect -4574 167818 -4338 168054
rect -4574 167498 -4338 167734
rect -4574 131818 -4338 132054
rect -4574 131498 -4338 131734
rect -4574 95818 -4338 96054
rect -4574 95498 -4338 95734
rect -4574 59818 -4338 60054
rect -4574 59498 -4338 59734
rect -4574 23818 -4338 24054
rect -4574 23498 -4338 23734
rect -3654 706442 -3418 706678
rect -3654 706122 -3418 706358
rect 4586 706442 4822 706678
rect 4586 706122 4822 706358
rect -3654 689818 -3418 690054
rect -3654 689498 -3418 689734
rect -3654 653818 -3418 654054
rect -3654 653498 -3418 653734
rect -3654 617818 -3418 618054
rect -3654 617498 -3418 617734
rect -3654 581818 -3418 582054
rect -3654 581498 -3418 581734
rect -3654 545818 -3418 546054
rect -3654 545498 -3418 545734
rect -3654 509818 -3418 510054
rect -3654 509498 -3418 509734
rect -3654 473818 -3418 474054
rect -3654 473498 -3418 473734
rect -3654 437818 -3418 438054
rect -3654 437498 -3418 437734
rect -3654 401818 -3418 402054
rect -3654 401498 -3418 401734
rect -3654 365818 -3418 366054
rect -3654 365498 -3418 365734
rect -3654 329818 -3418 330054
rect -3654 329498 -3418 329734
rect -3654 293818 -3418 294054
rect -3654 293498 -3418 293734
rect -3654 257818 -3418 258054
rect -3654 257498 -3418 257734
rect -3654 221818 -3418 222054
rect -3654 221498 -3418 221734
rect -3654 185818 -3418 186054
rect -3654 185498 -3418 185734
rect -3654 149818 -3418 150054
rect -3654 149498 -3418 149734
rect -3654 113818 -3418 114054
rect -3654 113498 -3418 113734
rect -3654 77818 -3418 78054
rect -3654 77498 -3418 77734
rect -3654 41818 -3418 42054
rect -3654 41498 -3418 41734
rect -3654 5818 -3418 6054
rect -3654 5498 -3418 5734
rect -2734 705522 -2498 705758
rect -2734 705202 -2498 705438
rect -2734 668218 -2498 668454
rect -2734 667898 -2498 668134
rect -2734 632218 -2498 632454
rect -2734 631898 -2498 632134
rect -2734 596218 -2498 596454
rect -2734 595898 -2498 596134
rect -2734 560218 -2498 560454
rect -2734 559898 -2498 560134
rect -2734 524218 -2498 524454
rect -2734 523898 -2498 524134
rect -2734 488218 -2498 488454
rect -2734 487898 -2498 488134
rect -2734 452218 -2498 452454
rect -2734 451898 -2498 452134
rect -2734 416218 -2498 416454
rect -2734 415898 -2498 416134
rect -2734 380218 -2498 380454
rect -2734 379898 -2498 380134
rect -2734 344218 -2498 344454
rect -2734 343898 -2498 344134
rect -2734 308218 -2498 308454
rect -2734 307898 -2498 308134
rect -2734 272218 -2498 272454
rect -2734 271898 -2498 272134
rect -2734 236218 -2498 236454
rect -2734 235898 -2498 236134
rect -2734 200218 -2498 200454
rect -2734 199898 -2498 200134
rect -2734 164218 -2498 164454
rect -2734 163898 -2498 164134
rect -2734 128218 -2498 128454
rect -2734 127898 -2498 128134
rect -2734 92218 -2498 92454
rect -2734 91898 -2498 92134
rect -2734 56218 -2498 56454
rect -2734 55898 -2498 56134
rect -2734 20218 -2498 20454
rect -2734 19898 -2498 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2734 -1502 -2498 -1266
rect -2734 -1822 -2498 -1586
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3654 -2422 -3418 -2186
rect -3654 -2742 -3418 -2506
rect 4586 -2422 4822 -2186
rect 4586 -2742 4822 -2506
rect -4574 -3342 -4338 -3106
rect -4574 -3662 -4338 -3426
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5494 -4262 -5258 -4026
rect -5494 -4582 -5258 -4346
rect 8186 -4262 8422 -4026
rect 8186 -4582 8422 -4346
rect -6414 -5182 -6178 -4946
rect -6414 -5502 -6178 -5266
rect 29786 711042 30022 711278
rect 29786 710722 30022 710958
rect 26186 709202 26422 709438
rect 26186 708882 26422 709118
rect 22586 707362 22822 707598
rect 22586 707042 22822 707278
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7334 -6102 -7098 -5866
rect -7334 -6422 -7098 -6186
rect 18986 705522 19222 705758
rect 18986 705202 19222 705438
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1502 19222 -1266
rect 18986 -1822 19222 -1586
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3342 22822 -3106
rect 22586 -3662 22822 -3426
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5182 26422 -4946
rect 26186 -5502 26422 -5266
rect 47786 710122 48022 710358
rect 47786 709802 48022 710038
rect 44186 708282 44422 708518
rect 44186 707962 44422 708198
rect 40586 706442 40822 706678
rect 40586 706122 40822 706358
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6102 12022 -5866
rect 11786 -6422 12022 -6186
rect -8254 -7022 -8018 -6786
rect -8254 -7342 -8018 -7106
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2422 40822 -2186
rect 40586 -2742 40822 -2506
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4262 44422 -4026
rect 44186 -4582 44422 -4346
rect 65786 711042 66022 711278
rect 65786 710722 66022 710958
rect 62186 709202 62422 709438
rect 62186 708882 62422 709118
rect 58586 707362 58822 707598
rect 58586 707042 58822 707278
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7022 30022 -6786
rect 29786 -7342 30022 -7106
rect 54986 705522 55222 705758
rect 54986 705202 55222 705438
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1502 55222 -1266
rect 54986 -1822 55222 -1586
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3342 58822 -3106
rect 58586 -3662 58822 -3426
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 62186 531418 62422 531654
rect 62186 531098 62422 531334
rect 62186 495418 62422 495654
rect 62186 495098 62422 495334
rect 62186 459418 62422 459654
rect 62186 459098 62422 459334
rect 62186 423418 62422 423654
rect 62186 423098 62422 423334
rect 62186 387418 62422 387654
rect 62186 387098 62422 387334
rect 62186 351418 62422 351654
rect 62186 351098 62422 351334
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5182 62422 -4946
rect 62186 -5502 62422 -5266
rect 83786 710122 84022 710358
rect 83786 709802 84022 710038
rect 80186 708282 80422 708518
rect 80186 707962 80422 708198
rect 76586 706442 76822 706678
rect 76586 706122 76822 706358
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 65786 535018 66022 535254
rect 65786 534698 66022 534934
rect 65786 499018 66022 499254
rect 65786 498698 66022 498934
rect 65786 463018 66022 463254
rect 65786 462698 66022 462934
rect 65786 427018 66022 427254
rect 65786 426698 66022 426934
rect 65786 391018 66022 391254
rect 65786 390698 66022 390934
rect 65786 355018 66022 355254
rect 65786 354698 66022 354934
rect 65786 319018 66022 319254
rect 65786 318698 66022 318934
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6102 48022 -5866
rect 47786 -6422 48022 -6186
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 76586 365818 76822 366054
rect 76586 365498 76822 365734
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2422 76822 -2186
rect 76586 -2742 76822 -2506
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 80186 621418 80422 621654
rect 80186 621098 80422 621334
rect 80186 585418 80422 585654
rect 80186 585098 80422 585334
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 80186 513418 80422 513654
rect 80186 513098 80422 513334
rect 80186 477418 80422 477654
rect 80186 477098 80422 477334
rect 80186 441418 80422 441654
rect 80186 441098 80422 441334
rect 80186 405418 80422 405654
rect 80186 405098 80422 405334
rect 80186 369418 80422 369654
rect 80186 369098 80422 369334
rect 80186 333418 80422 333654
rect 80186 333098 80422 333334
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4262 80422 -4026
rect 80186 -4582 80422 -4346
rect 101786 711042 102022 711278
rect 101786 710722 102022 710958
rect 98186 709202 98422 709438
rect 98186 708882 98422 709118
rect 94586 707362 94822 707598
rect 94586 707042 94822 707278
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 83786 625018 84022 625254
rect 83786 624698 84022 624934
rect 83786 589018 84022 589254
rect 83786 588698 84022 588934
rect 83786 553018 84022 553254
rect 83786 552698 84022 552934
rect 83786 517018 84022 517254
rect 83786 516698 84022 516934
rect 83786 481018 84022 481254
rect 83786 480698 84022 480934
rect 83786 445018 84022 445254
rect 83786 444698 84022 444934
rect 83786 409018 84022 409254
rect 83786 408698 84022 408934
rect 83786 373018 84022 373254
rect 83786 372698 84022 372934
rect 83786 337018 84022 337254
rect 83786 336698 84022 336934
rect 83786 301018 84022 301254
rect 83786 300698 84022 300934
rect 83786 265018 84022 265254
rect 83786 264698 84022 264934
rect 83786 229018 84022 229254
rect 83786 228698 84022 228934
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7022 66022 -6786
rect 65786 -7342 66022 -7106
rect 90986 705522 91222 705758
rect 90986 705202 91222 705438
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 90986 524218 91222 524454
rect 90986 523898 91222 524134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 90986 416218 91222 416454
rect 90986 415898 91222 416134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1502 91222 -1266
rect 90986 -1822 91222 -1586
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 94586 599818 94822 600054
rect 94586 599498 94822 599734
rect 94586 563818 94822 564054
rect 94586 563498 94822 563734
rect 94586 527818 94822 528054
rect 94586 527498 94822 527734
rect 94586 491818 94822 492054
rect 94586 491498 94822 491734
rect 94586 455818 94822 456054
rect 94586 455498 94822 455734
rect 94586 419818 94822 420054
rect 94586 419498 94822 419734
rect 94586 383818 94822 384054
rect 94586 383498 94822 383734
rect 94586 347818 94822 348054
rect 94586 347498 94822 347734
rect 94586 311818 94822 312054
rect 94586 311498 94822 311734
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3342 94822 -3106
rect 94586 -3662 94822 -3426
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 98186 639418 98422 639654
rect 98186 639098 98422 639334
rect 98186 603418 98422 603654
rect 98186 603098 98422 603334
rect 98186 567418 98422 567654
rect 98186 567098 98422 567334
rect 98186 531418 98422 531654
rect 98186 531098 98422 531334
rect 98186 495418 98422 495654
rect 98186 495098 98422 495334
rect 98186 459418 98422 459654
rect 98186 459098 98422 459334
rect 98186 423418 98422 423654
rect 98186 423098 98422 423334
rect 98186 387418 98422 387654
rect 98186 387098 98422 387334
rect 98186 351418 98422 351654
rect 98186 351098 98422 351334
rect 98186 315418 98422 315654
rect 98186 315098 98422 315334
rect 98186 279418 98422 279654
rect 98186 279098 98422 279334
rect 98186 243418 98422 243654
rect 98186 243098 98422 243334
rect 98186 207418 98422 207654
rect 98186 207098 98422 207334
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5182 98422 -4946
rect 98186 -5502 98422 -5266
rect 119786 710122 120022 710358
rect 119786 709802 120022 710038
rect 116186 708282 116422 708518
rect 116186 707962 116422 708198
rect 112586 706442 112822 706678
rect 112586 706122 112822 706358
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 101786 643018 102022 643254
rect 101786 642698 102022 642934
rect 101786 607018 102022 607254
rect 101786 606698 102022 606934
rect 101786 571018 102022 571254
rect 101786 570698 102022 570934
rect 101786 535018 102022 535254
rect 101786 534698 102022 534934
rect 101786 499018 102022 499254
rect 101786 498698 102022 498934
rect 101786 463018 102022 463254
rect 101786 462698 102022 462934
rect 101786 427018 102022 427254
rect 101786 426698 102022 426934
rect 101786 391018 102022 391254
rect 101786 390698 102022 390934
rect 101786 355018 102022 355254
rect 101786 354698 102022 354934
rect 101786 319018 102022 319254
rect 101786 318698 102022 318934
rect 101786 283018 102022 283254
rect 101786 282698 102022 282934
rect 101786 247018 102022 247254
rect 101786 246698 102022 246934
rect 101786 211018 102022 211254
rect 101786 210698 102022 210934
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6102 84022 -5866
rect 83786 -6422 84022 -6186
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 112586 581818 112822 582054
rect 112586 581498 112822 581734
rect 112586 545818 112822 546054
rect 112586 545498 112822 545734
rect 112586 509818 112822 510054
rect 112586 509498 112822 509734
rect 112586 473818 112822 474054
rect 112586 473498 112822 473734
rect 112586 437818 112822 438054
rect 112586 437498 112822 437734
rect 112586 401818 112822 402054
rect 112586 401498 112822 401734
rect 112586 365818 112822 366054
rect 112586 365498 112822 365734
rect 112586 329818 112822 330054
rect 112586 329498 112822 329734
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2422 112822 -2186
rect 112586 -2742 112822 -2506
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 116186 621418 116422 621654
rect 116186 621098 116422 621334
rect 116186 585418 116422 585654
rect 116186 585098 116422 585334
rect 116186 549418 116422 549654
rect 116186 549098 116422 549334
rect 116186 513418 116422 513654
rect 116186 513098 116422 513334
rect 116186 477418 116422 477654
rect 116186 477098 116422 477334
rect 116186 441418 116422 441654
rect 116186 441098 116422 441334
rect 116186 405418 116422 405654
rect 116186 405098 116422 405334
rect 116186 369418 116422 369654
rect 116186 369098 116422 369334
rect 116186 333418 116422 333654
rect 116186 333098 116422 333334
rect 116186 297418 116422 297654
rect 116186 297098 116422 297334
rect 116186 261418 116422 261654
rect 116186 261098 116422 261334
rect 116186 225418 116422 225654
rect 116186 225098 116422 225334
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4262 116422 -4026
rect 116186 -4582 116422 -4346
rect 137786 711042 138022 711278
rect 137786 710722 138022 710958
rect 134186 709202 134422 709438
rect 134186 708882 134422 709118
rect 130586 707362 130822 707598
rect 130586 707042 130822 707278
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 119786 625018 120022 625254
rect 119786 624698 120022 624934
rect 119786 589018 120022 589254
rect 119786 588698 120022 588934
rect 119786 553018 120022 553254
rect 119786 552698 120022 552934
rect 119786 517018 120022 517254
rect 119786 516698 120022 516934
rect 119786 481018 120022 481254
rect 119786 480698 120022 480934
rect 119786 445018 120022 445254
rect 119786 444698 120022 444934
rect 119786 409018 120022 409254
rect 119786 408698 120022 408934
rect 119786 373018 120022 373254
rect 119786 372698 120022 372934
rect 119786 337018 120022 337254
rect 119786 336698 120022 336934
rect 119786 301018 120022 301254
rect 119786 300698 120022 300934
rect 119786 265018 120022 265254
rect 119786 264698 120022 264934
rect 119786 229018 120022 229254
rect 119786 228698 120022 228934
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7022 102022 -6786
rect 101786 -7342 102022 -7106
rect 126986 705522 127222 705758
rect 126986 705202 127222 705438
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 126986 416218 127222 416454
rect 126986 415898 127222 416134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1502 127222 -1266
rect 126986 -1822 127222 -1586
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 130586 599818 130822 600054
rect 130586 599498 130822 599734
rect 130586 563818 130822 564054
rect 130586 563498 130822 563734
rect 130586 527818 130822 528054
rect 130586 527498 130822 527734
rect 130586 491818 130822 492054
rect 130586 491498 130822 491734
rect 130586 455818 130822 456054
rect 130586 455498 130822 455734
rect 130586 419818 130822 420054
rect 130586 419498 130822 419734
rect 130586 383818 130822 384054
rect 130586 383498 130822 383734
rect 130586 347818 130822 348054
rect 130586 347498 130822 347734
rect 130586 311818 130822 312054
rect 130586 311498 130822 311734
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3342 130822 -3106
rect 130586 -3662 130822 -3426
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 134186 639418 134422 639654
rect 134186 639098 134422 639334
rect 134186 603418 134422 603654
rect 134186 603098 134422 603334
rect 134186 567418 134422 567654
rect 134186 567098 134422 567334
rect 134186 531418 134422 531654
rect 134186 531098 134422 531334
rect 134186 495418 134422 495654
rect 134186 495098 134422 495334
rect 134186 459418 134422 459654
rect 134186 459098 134422 459334
rect 134186 423418 134422 423654
rect 134186 423098 134422 423334
rect 134186 387418 134422 387654
rect 134186 387098 134422 387334
rect 134186 351418 134422 351654
rect 134186 351098 134422 351334
rect 134186 315418 134422 315654
rect 134186 315098 134422 315334
rect 134186 279418 134422 279654
rect 134186 279098 134422 279334
rect 134186 243418 134422 243654
rect 134186 243098 134422 243334
rect 134186 207418 134422 207654
rect 134186 207098 134422 207334
rect 134186 171418 134422 171654
rect 134186 171098 134422 171334
rect 134186 135418 134422 135654
rect 134186 135098 134422 135334
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5182 134422 -4946
rect 134186 -5502 134422 -5266
rect 155786 710122 156022 710358
rect 155786 709802 156022 710038
rect 152186 708282 152422 708518
rect 152186 707962 152422 708198
rect 148586 706442 148822 706678
rect 148586 706122 148822 706358
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 137786 643018 138022 643254
rect 137786 642698 138022 642934
rect 137786 607018 138022 607254
rect 137786 606698 138022 606934
rect 137786 571018 138022 571254
rect 137786 570698 138022 570934
rect 137786 535018 138022 535254
rect 137786 534698 138022 534934
rect 137786 499018 138022 499254
rect 137786 498698 138022 498934
rect 137786 463018 138022 463254
rect 137786 462698 138022 462934
rect 137786 427018 138022 427254
rect 137786 426698 138022 426934
rect 137786 391018 138022 391254
rect 137786 390698 138022 390934
rect 137786 355018 138022 355254
rect 137786 354698 138022 354934
rect 137786 319018 138022 319254
rect 137786 318698 138022 318934
rect 137786 283018 138022 283254
rect 137786 282698 138022 282934
rect 137786 247018 138022 247254
rect 137786 246698 138022 246934
rect 137786 211018 138022 211254
rect 137786 210698 138022 210934
rect 137786 175018 138022 175254
rect 137786 174698 138022 174934
rect 137786 139018 138022 139254
rect 137786 138698 138022 138934
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6102 120022 -5866
rect 119786 -6422 120022 -6186
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 144986 506218 145222 506454
rect 144986 505898 145222 506134
rect 144986 470218 145222 470454
rect 144986 469898 145222 470134
rect 144986 434218 145222 434454
rect 144986 433898 145222 434134
rect 144986 398218 145222 398454
rect 144986 397898 145222 398134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 148586 509818 148822 510054
rect 148586 509498 148822 509734
rect 148586 473818 148822 474054
rect 148586 473498 148822 473734
rect 148586 437818 148822 438054
rect 148586 437498 148822 437734
rect 148586 401818 148822 402054
rect 148586 401498 148822 401734
rect 148586 365818 148822 366054
rect 148586 365498 148822 365734
rect 148586 329818 148822 330054
rect 148586 329498 148822 329734
rect 148586 293818 148822 294054
rect 148586 293498 148822 293734
rect 148586 257818 148822 258054
rect 148586 257498 148822 257734
rect 148586 221818 148822 222054
rect 148586 221498 148822 221734
rect 148586 185818 148822 186054
rect 148586 185498 148822 185734
rect 148586 149818 148822 150054
rect 148586 149498 148822 149734
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2422 148822 -2186
rect 148586 -2742 148822 -2506
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 152186 513418 152422 513654
rect 152186 513098 152422 513334
rect 152186 477418 152422 477654
rect 152186 477098 152422 477334
rect 152186 441418 152422 441654
rect 152186 441098 152422 441334
rect 152186 405418 152422 405654
rect 152186 405098 152422 405334
rect 152186 369418 152422 369654
rect 152186 369098 152422 369334
rect 152186 333418 152422 333654
rect 152186 333098 152422 333334
rect 152186 297418 152422 297654
rect 152186 297098 152422 297334
rect 152186 261418 152422 261654
rect 152186 261098 152422 261334
rect 152186 225418 152422 225654
rect 152186 225098 152422 225334
rect 152186 189418 152422 189654
rect 152186 189098 152422 189334
rect 152186 153418 152422 153654
rect 152186 153098 152422 153334
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4262 152422 -4026
rect 152186 -4582 152422 -4346
rect 173786 711042 174022 711278
rect 173786 710722 174022 710958
rect 170186 709202 170422 709438
rect 170186 708882 170422 709118
rect 166586 707362 166822 707598
rect 166586 707042 166822 707278
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 155786 517018 156022 517254
rect 155786 516698 156022 516934
rect 155786 481018 156022 481254
rect 155786 480698 156022 480934
rect 155786 445018 156022 445254
rect 155786 444698 156022 444934
rect 155786 409018 156022 409254
rect 155786 408698 156022 408934
rect 155786 373018 156022 373254
rect 155786 372698 156022 372934
rect 155786 337018 156022 337254
rect 155786 336698 156022 336934
rect 155786 301018 156022 301254
rect 155786 300698 156022 300934
rect 155786 265018 156022 265254
rect 155786 264698 156022 264934
rect 155786 229018 156022 229254
rect 155786 228698 156022 228934
rect 155786 193018 156022 193254
rect 155786 192698 156022 192934
rect 155786 157018 156022 157254
rect 155786 156698 156022 156934
rect 155786 121018 156022 121254
rect 155786 120698 156022 120934
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7022 138022 -6786
rect 137786 -7342 138022 -7106
rect 162986 705522 163222 705758
rect 162986 705202 163222 705438
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 162986 416218 163222 416454
rect 162986 415898 163222 416134
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 162986 344218 163222 344454
rect 162986 343898 163222 344134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 162986 200218 163222 200454
rect 162986 199898 163222 200134
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1502 163222 -1266
rect 162986 -1822 163222 -1586
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 166586 527818 166822 528054
rect 166586 527498 166822 527734
rect 166586 491818 166822 492054
rect 166586 491498 166822 491734
rect 166586 455818 166822 456054
rect 166586 455498 166822 455734
rect 166586 419818 166822 420054
rect 166586 419498 166822 419734
rect 166586 383818 166822 384054
rect 166586 383498 166822 383734
rect 166586 347818 166822 348054
rect 166586 347498 166822 347734
rect 166586 311818 166822 312054
rect 166586 311498 166822 311734
rect 166586 275818 166822 276054
rect 166586 275498 166822 275734
rect 166586 239818 166822 240054
rect 166586 239498 166822 239734
rect 166586 203818 166822 204054
rect 166586 203498 166822 203734
rect 166586 167818 166822 168054
rect 166586 167498 166822 167734
rect 166586 131818 166822 132054
rect 166586 131498 166822 131734
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3342 166822 -3106
rect 166586 -3662 166822 -3426
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 170186 531418 170422 531654
rect 170186 531098 170422 531334
rect 170186 495418 170422 495654
rect 170186 495098 170422 495334
rect 170186 459418 170422 459654
rect 170186 459098 170422 459334
rect 170186 423418 170422 423654
rect 170186 423098 170422 423334
rect 170186 387418 170422 387654
rect 170186 387098 170422 387334
rect 170186 351418 170422 351654
rect 170186 351098 170422 351334
rect 170186 315418 170422 315654
rect 170186 315098 170422 315334
rect 170186 279418 170422 279654
rect 170186 279098 170422 279334
rect 170186 243418 170422 243654
rect 170186 243098 170422 243334
rect 170186 207418 170422 207654
rect 170186 207098 170422 207334
rect 170186 171418 170422 171654
rect 170186 171098 170422 171334
rect 170186 135418 170422 135654
rect 170186 135098 170422 135334
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5182 170422 -4946
rect 170186 -5502 170422 -5266
rect 191786 710122 192022 710358
rect 191786 709802 192022 710038
rect 188186 708282 188422 708518
rect 188186 707962 188422 708198
rect 184586 706442 184822 706678
rect 184586 706122 184822 706358
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 173786 535018 174022 535254
rect 173786 534698 174022 534934
rect 173786 499018 174022 499254
rect 173786 498698 174022 498934
rect 173786 463018 174022 463254
rect 173786 462698 174022 462934
rect 173786 427018 174022 427254
rect 173786 426698 174022 426934
rect 173786 391018 174022 391254
rect 173786 390698 174022 390934
rect 173786 355018 174022 355254
rect 173786 354698 174022 354934
rect 173786 319018 174022 319254
rect 173786 318698 174022 318934
rect 173786 283018 174022 283254
rect 173786 282698 174022 282934
rect 173786 247018 174022 247254
rect 173786 246698 174022 246934
rect 173786 211018 174022 211254
rect 173786 210698 174022 210934
rect 173786 175018 174022 175254
rect 173786 174698 174022 174934
rect 173786 139018 174022 139254
rect 173786 138698 174022 138934
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6102 156022 -5866
rect 155786 -6422 156022 -6186
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 180986 506218 181222 506454
rect 180986 505898 181222 506134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 180986 434218 181222 434454
rect 180986 433898 181222 434134
rect 180986 398218 181222 398454
rect 180986 397898 181222 398134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 180986 326218 181222 326454
rect 180986 325898 181222 326134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 180986 218218 181222 218454
rect 180986 217898 181222 218134
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 184586 509818 184822 510054
rect 184586 509498 184822 509734
rect 184586 473818 184822 474054
rect 184586 473498 184822 473734
rect 184586 437818 184822 438054
rect 184586 437498 184822 437734
rect 184586 401818 184822 402054
rect 184586 401498 184822 401734
rect 184586 365818 184822 366054
rect 184586 365498 184822 365734
rect 184586 329818 184822 330054
rect 184586 329498 184822 329734
rect 184586 293818 184822 294054
rect 184586 293498 184822 293734
rect 184586 257818 184822 258054
rect 184586 257498 184822 257734
rect 184586 221818 184822 222054
rect 184586 221498 184822 221734
rect 184586 185818 184822 186054
rect 184586 185498 184822 185734
rect 184586 149818 184822 150054
rect 184586 149498 184822 149734
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2422 184822 -2186
rect 184586 -2742 184822 -2506
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 188186 585418 188422 585654
rect 188186 585098 188422 585334
rect 188186 549418 188422 549654
rect 188186 549098 188422 549334
rect 188186 513418 188422 513654
rect 188186 513098 188422 513334
rect 188186 477418 188422 477654
rect 188186 477098 188422 477334
rect 188186 441418 188422 441654
rect 188186 441098 188422 441334
rect 188186 405418 188422 405654
rect 188186 405098 188422 405334
rect 188186 369418 188422 369654
rect 188186 369098 188422 369334
rect 188186 333418 188422 333654
rect 188186 333098 188422 333334
rect 188186 297418 188422 297654
rect 188186 297098 188422 297334
rect 188186 261418 188422 261654
rect 188186 261098 188422 261334
rect 188186 225418 188422 225654
rect 188186 225098 188422 225334
rect 188186 189418 188422 189654
rect 188186 189098 188422 189334
rect 188186 153418 188422 153654
rect 188186 153098 188422 153334
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4262 188422 -4026
rect 188186 -4582 188422 -4346
rect 209786 711042 210022 711278
rect 209786 710722 210022 710958
rect 206186 709202 206422 709438
rect 206186 708882 206422 709118
rect 202586 707362 202822 707598
rect 202586 707042 202822 707278
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 191786 625018 192022 625254
rect 191786 624698 192022 624934
rect 191786 589018 192022 589254
rect 191786 588698 192022 588934
rect 191786 553018 192022 553254
rect 191786 552698 192022 552934
rect 191786 517018 192022 517254
rect 191786 516698 192022 516934
rect 191786 481018 192022 481254
rect 191786 480698 192022 480934
rect 191786 445018 192022 445254
rect 191786 444698 192022 444934
rect 191786 409018 192022 409254
rect 191786 408698 192022 408934
rect 191786 373018 192022 373254
rect 191786 372698 192022 372934
rect 191786 337018 192022 337254
rect 191786 336698 192022 336934
rect 191786 301018 192022 301254
rect 191786 300698 192022 300934
rect 191786 265018 192022 265254
rect 191786 264698 192022 264934
rect 191786 229018 192022 229254
rect 191786 228698 192022 228934
rect 191786 193018 192022 193254
rect 191786 192698 192022 192934
rect 191786 157018 192022 157254
rect 191786 156698 192022 156934
rect 191786 121018 192022 121254
rect 191786 120698 192022 120934
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7022 174022 -6786
rect 173786 -7342 174022 -7106
rect 198986 705522 199222 705758
rect 198986 705202 199222 705438
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 198986 524218 199222 524454
rect 198986 523898 199222 524134
rect 198986 488218 199222 488454
rect 198986 487898 199222 488134
rect 198986 452218 199222 452454
rect 198986 451898 199222 452134
rect 198986 416218 199222 416454
rect 198986 415898 199222 416134
rect 198986 380218 199222 380454
rect 198986 379898 199222 380134
rect 198986 344218 199222 344454
rect 198986 343898 199222 344134
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 198986 272218 199222 272454
rect 198986 271898 199222 272134
rect 198986 236218 199222 236454
rect 198986 235898 199222 236134
rect 198986 200218 199222 200454
rect 198986 199898 199222 200134
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1502 199222 -1266
rect 198986 -1822 199222 -1586
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 202586 599818 202822 600054
rect 202586 599498 202822 599734
rect 202586 563818 202822 564054
rect 202586 563498 202822 563734
rect 202586 527818 202822 528054
rect 202586 527498 202822 527734
rect 202586 491818 202822 492054
rect 202586 491498 202822 491734
rect 202586 455818 202822 456054
rect 202586 455498 202822 455734
rect 202586 419818 202822 420054
rect 202586 419498 202822 419734
rect 202586 383818 202822 384054
rect 202586 383498 202822 383734
rect 202586 347818 202822 348054
rect 202586 347498 202822 347734
rect 202586 311818 202822 312054
rect 202586 311498 202822 311734
rect 202586 275818 202822 276054
rect 202586 275498 202822 275734
rect 202586 239818 202822 240054
rect 202586 239498 202822 239734
rect 202586 203818 202822 204054
rect 202586 203498 202822 203734
rect 202586 167818 202822 168054
rect 202586 167498 202822 167734
rect 202586 131818 202822 132054
rect 202586 131498 202822 131734
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3342 202822 -3106
rect 202586 -3662 202822 -3426
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 206186 639418 206422 639654
rect 206186 639098 206422 639334
rect 206186 603418 206422 603654
rect 206186 603098 206422 603334
rect 206186 567418 206422 567654
rect 206186 567098 206422 567334
rect 206186 531418 206422 531654
rect 206186 531098 206422 531334
rect 206186 495418 206422 495654
rect 206186 495098 206422 495334
rect 206186 459418 206422 459654
rect 206186 459098 206422 459334
rect 206186 423418 206422 423654
rect 206186 423098 206422 423334
rect 206186 387418 206422 387654
rect 206186 387098 206422 387334
rect 206186 351418 206422 351654
rect 206186 351098 206422 351334
rect 206186 315418 206422 315654
rect 206186 315098 206422 315334
rect 206186 279418 206422 279654
rect 206186 279098 206422 279334
rect 206186 243418 206422 243654
rect 206186 243098 206422 243334
rect 206186 207418 206422 207654
rect 206186 207098 206422 207334
rect 206186 171418 206422 171654
rect 206186 171098 206422 171334
rect 206186 135418 206422 135654
rect 206186 135098 206422 135334
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5182 206422 -4946
rect 206186 -5502 206422 -5266
rect 227786 710122 228022 710358
rect 227786 709802 228022 710038
rect 224186 708282 224422 708518
rect 224186 707962 224422 708198
rect 220586 706442 220822 706678
rect 220586 706122 220822 706358
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 209786 643018 210022 643254
rect 209786 642698 210022 642934
rect 209786 607018 210022 607254
rect 209786 606698 210022 606934
rect 209786 571018 210022 571254
rect 209786 570698 210022 570934
rect 209786 535018 210022 535254
rect 209786 534698 210022 534934
rect 209786 499018 210022 499254
rect 209786 498698 210022 498934
rect 209786 463018 210022 463254
rect 209786 462698 210022 462934
rect 209786 427018 210022 427254
rect 209786 426698 210022 426934
rect 209786 391018 210022 391254
rect 209786 390698 210022 390934
rect 209786 355018 210022 355254
rect 209786 354698 210022 354934
rect 209786 319018 210022 319254
rect 209786 318698 210022 318934
rect 209786 283018 210022 283254
rect 209786 282698 210022 282934
rect 209786 247018 210022 247254
rect 209786 246698 210022 246934
rect 209786 211018 210022 211254
rect 209786 210698 210022 210934
rect 209786 175018 210022 175254
rect 209786 174698 210022 174934
rect 209786 139018 210022 139254
rect 209786 138698 210022 138934
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6102 192022 -5866
rect 191786 -6422 192022 -6186
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 216986 542218 217222 542454
rect 216986 541898 217222 542134
rect 216986 506218 217222 506454
rect 216986 505898 217222 506134
rect 216986 470218 217222 470454
rect 216986 469898 217222 470134
rect 216986 434218 217222 434454
rect 216986 433898 217222 434134
rect 216986 398218 217222 398454
rect 216986 397898 217222 398134
rect 216986 362218 217222 362454
rect 216986 361898 217222 362134
rect 216986 326218 217222 326454
rect 216986 325898 217222 326134
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 216986 254218 217222 254454
rect 216986 253898 217222 254134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 220586 581818 220822 582054
rect 220586 581498 220822 581734
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 220586 509818 220822 510054
rect 220586 509498 220822 509734
rect 220586 473818 220822 474054
rect 220586 473498 220822 473734
rect 220586 437818 220822 438054
rect 220586 437498 220822 437734
rect 220586 401818 220822 402054
rect 220586 401498 220822 401734
rect 220586 365818 220822 366054
rect 220586 365498 220822 365734
rect 220586 329818 220822 330054
rect 220586 329498 220822 329734
rect 220586 293818 220822 294054
rect 220586 293498 220822 293734
rect 220586 257818 220822 258054
rect 220586 257498 220822 257734
rect 220586 221818 220822 222054
rect 220586 221498 220822 221734
rect 220586 185818 220822 186054
rect 220586 185498 220822 185734
rect 220586 149818 220822 150054
rect 220586 149498 220822 149734
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2422 220822 -2186
rect 220586 -2742 220822 -2506
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 224186 621418 224422 621654
rect 224186 621098 224422 621334
rect 224186 585418 224422 585654
rect 224186 585098 224422 585334
rect 224186 549418 224422 549654
rect 224186 549098 224422 549334
rect 224186 513418 224422 513654
rect 224186 513098 224422 513334
rect 224186 477418 224422 477654
rect 224186 477098 224422 477334
rect 224186 441418 224422 441654
rect 224186 441098 224422 441334
rect 224186 405418 224422 405654
rect 224186 405098 224422 405334
rect 224186 369418 224422 369654
rect 224186 369098 224422 369334
rect 224186 333418 224422 333654
rect 224186 333098 224422 333334
rect 224186 297418 224422 297654
rect 224186 297098 224422 297334
rect 224186 261418 224422 261654
rect 224186 261098 224422 261334
rect 224186 225418 224422 225654
rect 224186 225098 224422 225334
rect 224186 189418 224422 189654
rect 224186 189098 224422 189334
rect 224186 153418 224422 153654
rect 224186 153098 224422 153334
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4262 224422 -4026
rect 224186 -4582 224422 -4346
rect 245786 711042 246022 711278
rect 245786 710722 246022 710958
rect 242186 709202 242422 709438
rect 242186 708882 242422 709118
rect 238586 707362 238822 707598
rect 238586 707042 238822 707278
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 227786 625018 228022 625254
rect 227786 624698 228022 624934
rect 227786 589018 228022 589254
rect 227786 588698 228022 588934
rect 227786 553018 228022 553254
rect 227786 552698 228022 552934
rect 227786 517018 228022 517254
rect 227786 516698 228022 516934
rect 227786 481018 228022 481254
rect 227786 480698 228022 480934
rect 234986 705522 235222 705758
rect 234986 705202 235222 705438
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 234986 524218 235222 524454
rect 234986 523898 235222 524134
rect 234986 488218 235222 488454
rect 234986 487898 235222 488134
rect 227786 445018 228022 445254
rect 227786 444698 228022 444934
rect 227786 409018 228022 409254
rect 227786 408698 228022 408934
rect 227786 373018 228022 373254
rect 227786 372698 228022 372934
rect 227786 337018 228022 337254
rect 227786 336698 228022 336934
rect 227786 301018 228022 301254
rect 227786 300698 228022 300934
rect 227786 265018 228022 265254
rect 227786 264698 228022 264934
rect 227786 229018 228022 229254
rect 227786 228698 228022 228934
rect 227786 193018 228022 193254
rect 227786 192698 228022 192934
rect 227786 157018 228022 157254
rect 227786 156698 228022 156934
rect 227786 121018 228022 121254
rect 227786 120698 228022 120934
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 234986 452218 235222 452454
rect 234986 451898 235222 452134
rect 234986 416218 235222 416454
rect 234986 415898 235222 416134
rect 234986 380218 235222 380454
rect 234986 379898 235222 380134
rect 234986 344218 235222 344454
rect 234986 343898 235222 344134
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 234986 272218 235222 272454
rect 234986 271898 235222 272134
rect 234986 236218 235222 236454
rect 234986 235898 235222 236134
rect 234986 200218 235222 200454
rect 234986 199898 235222 200134
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7022 210022 -6786
rect 209786 -7342 210022 -7106
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 238586 599818 238822 600054
rect 238586 599498 238822 599734
rect 238586 563818 238822 564054
rect 238586 563498 238822 563734
rect 238586 527818 238822 528054
rect 238586 527498 238822 527734
rect 238586 491818 238822 492054
rect 238586 491498 238822 491734
rect 238586 455818 238822 456054
rect 238586 455498 238822 455734
rect 238586 419818 238822 420054
rect 238586 419498 238822 419734
rect 238586 383818 238822 384054
rect 238586 383498 238822 383734
rect 238586 347818 238822 348054
rect 238586 347498 238822 347734
rect 238586 311818 238822 312054
rect 238586 311498 238822 311734
rect 238586 275818 238822 276054
rect 238586 275498 238822 275734
rect 238586 239818 238822 240054
rect 238586 239498 238822 239734
rect 238586 203818 238822 204054
rect 238586 203498 238822 203734
rect 238586 167818 238822 168054
rect 238586 167498 238822 167734
rect 238586 131818 238822 132054
rect 238586 131498 238822 131734
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1502 235222 -1266
rect 234986 -1822 235222 -1586
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 242186 639418 242422 639654
rect 242186 639098 242422 639334
rect 242186 603418 242422 603654
rect 242186 603098 242422 603334
rect 242186 567418 242422 567654
rect 242186 567098 242422 567334
rect 242186 531418 242422 531654
rect 242186 531098 242422 531334
rect 242186 495418 242422 495654
rect 242186 495098 242422 495334
rect 242186 459418 242422 459654
rect 242186 459098 242422 459334
rect 242186 423418 242422 423654
rect 242186 423098 242422 423334
rect 242186 387418 242422 387654
rect 242186 387098 242422 387334
rect 242186 351418 242422 351654
rect 242186 351098 242422 351334
rect 242186 315418 242422 315654
rect 242186 315098 242422 315334
rect 242186 279418 242422 279654
rect 242186 279098 242422 279334
rect 242186 243418 242422 243654
rect 242186 243098 242422 243334
rect 242186 207418 242422 207654
rect 242186 207098 242422 207334
rect 242186 171418 242422 171654
rect 242186 171098 242422 171334
rect 263786 710122 264022 710358
rect 263786 709802 264022 710038
rect 260186 708282 260422 708518
rect 260186 707962 260422 708198
rect 256586 706442 256822 706678
rect 256586 706122 256822 706358
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 245786 643018 246022 643254
rect 245786 642698 246022 642934
rect 245786 607018 246022 607254
rect 245786 606698 246022 606934
rect 245786 571018 246022 571254
rect 245786 570698 246022 570934
rect 245786 535018 246022 535254
rect 245786 534698 246022 534934
rect 245786 499018 246022 499254
rect 245786 498698 246022 498934
rect 245786 463018 246022 463254
rect 245786 462698 246022 462934
rect 245786 427018 246022 427254
rect 245786 426698 246022 426934
rect 245786 391018 246022 391254
rect 245786 390698 246022 390934
rect 245786 355018 246022 355254
rect 245786 354698 246022 354934
rect 245786 319018 246022 319254
rect 245786 318698 246022 318934
rect 245786 283018 246022 283254
rect 245786 282698 246022 282934
rect 245786 247018 246022 247254
rect 245786 246698 246022 246934
rect 245786 211018 246022 211254
rect 245786 210698 246022 210934
rect 245786 175018 246022 175254
rect 245786 174698 246022 174934
rect 245786 139018 246022 139254
rect 245786 138698 246022 138934
rect 242186 135418 242422 135654
rect 242186 135098 242422 135334
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3342 238822 -3106
rect 238586 -3662 238822 -3426
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5182 242422 -4946
rect 242186 -5502 242422 -5266
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6102 228022 -5866
rect 227786 -6422 228022 -6186
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 252986 506218 253222 506454
rect 252986 505898 253222 506134
rect 252986 470218 253222 470454
rect 252986 469898 253222 470134
rect 252986 434218 253222 434454
rect 252986 433898 253222 434134
rect 252986 398218 253222 398454
rect 252986 397898 253222 398134
rect 252986 362218 253222 362454
rect 252986 361898 253222 362134
rect 252986 326218 253222 326454
rect 252986 325898 253222 326134
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 252986 254218 253222 254454
rect 252986 253898 253222 254134
rect 252986 218218 253222 218454
rect 252986 217898 253222 218134
rect 252986 182218 253222 182454
rect 252986 181898 253222 182134
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 256586 581818 256822 582054
rect 256586 581498 256822 581734
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 256586 509818 256822 510054
rect 256586 509498 256822 509734
rect 256586 473818 256822 474054
rect 256586 473498 256822 473734
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 260186 621418 260422 621654
rect 260186 621098 260422 621334
rect 260186 585418 260422 585654
rect 260186 585098 260422 585334
rect 260186 549418 260422 549654
rect 260186 549098 260422 549334
rect 260186 513418 260422 513654
rect 260186 513098 260422 513334
rect 260186 477418 260422 477654
rect 260186 477098 260422 477334
rect 256586 437818 256822 438054
rect 256586 437498 256822 437734
rect 256586 401818 256822 402054
rect 256586 401498 256822 401734
rect 256586 365818 256822 366054
rect 256586 365498 256822 365734
rect 256586 329818 256822 330054
rect 256586 329498 256822 329734
rect 256586 293818 256822 294054
rect 256586 293498 256822 293734
rect 256586 257818 256822 258054
rect 256586 257498 256822 257734
rect 256586 221818 256822 222054
rect 256586 221498 256822 221734
rect 256586 185818 256822 186054
rect 256586 185498 256822 185734
rect 256586 149818 256822 150054
rect 256586 149498 256822 149734
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 260186 441418 260422 441654
rect 260186 441098 260422 441334
rect 260186 405418 260422 405654
rect 260186 405098 260422 405334
rect 260186 369418 260422 369654
rect 260186 369098 260422 369334
rect 260186 333418 260422 333654
rect 260186 333098 260422 333334
rect 260186 297418 260422 297654
rect 260186 297098 260422 297334
rect 260186 261418 260422 261654
rect 260186 261098 260422 261334
rect 260186 225418 260422 225654
rect 260186 225098 260422 225334
rect 260186 189418 260422 189654
rect 260186 189098 260422 189334
rect 260186 153418 260422 153654
rect 260186 153098 260422 153334
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2422 256822 -2186
rect 256586 -2742 256822 -2506
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4262 260422 -4026
rect 260186 -4582 260422 -4346
rect 281786 711042 282022 711278
rect 281786 710722 282022 710958
rect 278186 709202 278422 709438
rect 278186 708882 278422 709118
rect 274586 707362 274822 707598
rect 274586 707042 274822 707278
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 263786 625018 264022 625254
rect 263786 624698 264022 624934
rect 263786 589018 264022 589254
rect 263786 588698 264022 588934
rect 263786 553018 264022 553254
rect 263786 552698 264022 552934
rect 263786 517018 264022 517254
rect 263786 516698 264022 516934
rect 263786 481018 264022 481254
rect 263786 480698 264022 480934
rect 263786 445018 264022 445254
rect 263786 444698 264022 444934
rect 263786 409018 264022 409254
rect 263786 408698 264022 408934
rect 263786 373018 264022 373254
rect 263786 372698 264022 372934
rect 270986 705522 271222 705758
rect 270986 705202 271222 705438
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 270986 416218 271222 416454
rect 270986 415898 271222 416134
rect 270986 380218 271222 380454
rect 270986 379898 271222 380134
rect 270986 344218 271222 344454
rect 270986 343898 271222 344134
rect 263786 337018 264022 337254
rect 263786 336698 264022 336934
rect 263786 301018 264022 301254
rect 263786 300698 264022 300934
rect 263786 265018 264022 265254
rect 263786 264698 264022 264934
rect 263786 229018 264022 229254
rect 263786 228698 264022 228934
rect 263786 193018 264022 193254
rect 263786 192698 264022 192934
rect 263786 157018 264022 157254
rect 263786 156698 264022 156934
rect 263786 121018 264022 121254
rect 263786 120698 264022 120934
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7022 246022 -6786
rect 245786 -7342 246022 -7106
rect 270986 -1502 271222 -1266
rect 270986 -1822 271222 -1586
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 274586 527818 274822 528054
rect 274586 527498 274822 527734
rect 274586 491818 274822 492054
rect 274586 491498 274822 491734
rect 274586 455818 274822 456054
rect 274586 455498 274822 455734
rect 274586 419818 274822 420054
rect 274586 419498 274822 419734
rect 274586 383818 274822 384054
rect 274586 383498 274822 383734
rect 274586 347818 274822 348054
rect 274586 347498 274822 347734
rect 274586 311818 274822 312054
rect 274586 311498 274822 311734
rect 274586 275818 274822 276054
rect 274586 275498 274822 275734
rect 274586 239818 274822 240054
rect 274586 239498 274822 239734
rect 274586 203818 274822 204054
rect 274586 203498 274822 203734
rect 274586 167818 274822 168054
rect 274586 167498 274822 167734
rect 274586 131818 274822 132054
rect 274586 131498 274822 131734
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 278186 531418 278422 531654
rect 278186 531098 278422 531334
rect 278186 495418 278422 495654
rect 278186 495098 278422 495334
rect 278186 459418 278422 459654
rect 278186 459098 278422 459334
rect 278186 423418 278422 423654
rect 278186 423098 278422 423334
rect 278186 387418 278422 387654
rect 278186 387098 278422 387334
rect 278186 351418 278422 351654
rect 278186 351098 278422 351334
rect 278186 315418 278422 315654
rect 278186 315098 278422 315334
rect 278186 279418 278422 279654
rect 278186 279098 278422 279334
rect 278186 243418 278422 243654
rect 278186 243098 278422 243334
rect 278186 207418 278422 207654
rect 278186 207098 278422 207334
rect 278186 171418 278422 171654
rect 278186 171098 278422 171334
rect 278186 135418 278422 135654
rect 278186 135098 278422 135334
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 278186 63098 278422 63334
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3342 274822 -3106
rect 274586 -3662 274822 -3426
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5182 278422 -4946
rect 278186 -5502 278422 -5266
rect 299786 710122 300022 710358
rect 299786 709802 300022 710038
rect 296186 708282 296422 708518
rect 296186 707962 296422 708198
rect 292586 706442 292822 706678
rect 292586 706122 292822 706358
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 281786 535018 282022 535254
rect 281786 534698 282022 534934
rect 281786 499018 282022 499254
rect 281786 498698 282022 498934
rect 281786 463018 282022 463254
rect 281786 462698 282022 462934
rect 281786 427018 282022 427254
rect 281786 426698 282022 426934
rect 281786 391018 282022 391254
rect 281786 390698 282022 390934
rect 281786 355018 282022 355254
rect 281786 354698 282022 354934
rect 281786 319018 282022 319254
rect 281786 318698 282022 318934
rect 281786 283018 282022 283254
rect 281786 282698 282022 282934
rect 281786 247018 282022 247254
rect 281786 246698 282022 246934
rect 281786 211018 282022 211254
rect 281786 210698 282022 210934
rect 281786 175018 282022 175254
rect 281786 174698 282022 174934
rect 281786 139018 282022 139254
rect 281786 138698 282022 138934
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6102 264022 -5866
rect 263786 -6422 264022 -6186
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 288986 326218 289222 326454
rect 288986 325898 289222 326134
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 292586 473818 292822 474054
rect 292586 473498 292822 473734
rect 292586 437818 292822 438054
rect 292586 437498 292822 437734
rect 292586 401818 292822 402054
rect 292586 401498 292822 401734
rect 292586 365818 292822 366054
rect 292586 365498 292822 365734
rect 292586 329818 292822 330054
rect 292586 329498 292822 329734
rect 292586 293818 292822 294054
rect 292586 293498 292822 293734
rect 292586 257818 292822 258054
rect 292586 257498 292822 257734
rect 292586 221818 292822 222054
rect 292586 221498 292822 221734
rect 292586 185818 292822 186054
rect 292586 185498 292822 185734
rect 292586 149818 292822 150054
rect 292586 149498 292822 149734
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2422 292822 -2186
rect 292586 -2742 292822 -2506
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 296186 513418 296422 513654
rect 296186 513098 296422 513334
rect 296186 477418 296422 477654
rect 296186 477098 296422 477334
rect 296186 441418 296422 441654
rect 296186 441098 296422 441334
rect 296186 405418 296422 405654
rect 296186 405098 296422 405334
rect 296186 369418 296422 369654
rect 296186 369098 296422 369334
rect 296186 333418 296422 333654
rect 296186 333098 296422 333334
rect 296186 297418 296422 297654
rect 296186 297098 296422 297334
rect 296186 261418 296422 261654
rect 296186 261098 296422 261334
rect 296186 225418 296422 225654
rect 296186 225098 296422 225334
rect 296186 189418 296422 189654
rect 296186 189098 296422 189334
rect 296186 153418 296422 153654
rect 296186 153098 296422 153334
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4262 296422 -4026
rect 296186 -4582 296422 -4346
rect 317786 711042 318022 711278
rect 317786 710722 318022 710958
rect 314186 709202 314422 709438
rect 314186 708882 314422 709118
rect 310586 707362 310822 707598
rect 310586 707042 310822 707278
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 299786 589018 300022 589254
rect 299786 588698 300022 588934
rect 299786 553018 300022 553254
rect 299786 552698 300022 552934
rect 299786 517018 300022 517254
rect 299786 516698 300022 516934
rect 299786 481018 300022 481254
rect 299786 480698 300022 480934
rect 299786 445018 300022 445254
rect 299786 444698 300022 444934
rect 299786 409018 300022 409254
rect 299786 408698 300022 408934
rect 299786 373018 300022 373254
rect 299786 372698 300022 372934
rect 299786 337018 300022 337254
rect 299786 336698 300022 336934
rect 299786 301018 300022 301254
rect 299786 300698 300022 300934
rect 299786 265018 300022 265254
rect 299786 264698 300022 264934
rect 299786 229018 300022 229254
rect 299786 228698 300022 228934
rect 299786 193018 300022 193254
rect 299786 192698 300022 192934
rect 299786 157018 300022 157254
rect 299786 156698 300022 156934
rect 299786 121018 300022 121254
rect 299786 120698 300022 120934
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 306986 705522 307222 705758
rect 306986 705202 307222 705438
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 306986 344218 307222 344454
rect 306986 343898 307222 344134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 306986 200218 307222 200454
rect 306986 199898 307222 200134
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7022 282022 -6786
rect 281786 -7342 282022 -7106
rect 306986 -1502 307222 -1266
rect 306986 -1822 307222 -1586
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 310586 599818 310822 600054
rect 310586 599498 310822 599734
rect 310586 563818 310822 564054
rect 310586 563498 310822 563734
rect 310586 527818 310822 528054
rect 310586 527498 310822 527734
rect 310586 491818 310822 492054
rect 310586 491498 310822 491734
rect 310586 455818 310822 456054
rect 310586 455498 310822 455734
rect 310586 419818 310822 420054
rect 310586 419498 310822 419734
rect 310586 383818 310822 384054
rect 310586 383498 310822 383734
rect 310586 347818 310822 348054
rect 310586 347498 310822 347734
rect 310586 311818 310822 312054
rect 310586 311498 310822 311734
rect 310586 275818 310822 276054
rect 310586 275498 310822 275734
rect 310586 239818 310822 240054
rect 310586 239498 310822 239734
rect 310586 203818 310822 204054
rect 310586 203498 310822 203734
rect 310586 167818 310822 168054
rect 310586 167498 310822 167734
rect 310586 131818 310822 132054
rect 310586 131498 310822 131734
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 314186 603418 314422 603654
rect 314186 603098 314422 603334
rect 314186 567418 314422 567654
rect 314186 567098 314422 567334
rect 314186 531418 314422 531654
rect 314186 531098 314422 531334
rect 314186 495418 314422 495654
rect 314186 495098 314422 495334
rect 314186 459418 314422 459654
rect 314186 459098 314422 459334
rect 314186 423418 314422 423654
rect 314186 423098 314422 423334
rect 314186 387418 314422 387654
rect 314186 387098 314422 387334
rect 314186 351418 314422 351654
rect 314186 351098 314422 351334
rect 314186 315418 314422 315654
rect 314186 315098 314422 315334
rect 314186 279418 314422 279654
rect 314186 279098 314422 279334
rect 314186 243418 314422 243654
rect 314186 243098 314422 243334
rect 314186 207418 314422 207654
rect 314186 207098 314422 207334
rect 314186 171418 314422 171654
rect 314186 171098 314422 171334
rect 314186 135418 314422 135654
rect 314186 135098 314422 135334
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 335786 710122 336022 710358
rect 335786 709802 336022 710038
rect 332186 708282 332422 708518
rect 332186 707962 332422 708198
rect 328586 706442 328822 706678
rect 328586 706122 328822 706358
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 317786 607018 318022 607254
rect 317786 606698 318022 606934
rect 317786 571018 318022 571254
rect 317786 570698 318022 570934
rect 317786 535018 318022 535254
rect 317786 534698 318022 534934
rect 317786 499018 318022 499254
rect 317786 498698 318022 498934
rect 317786 463018 318022 463254
rect 317786 462698 318022 462934
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 324986 578218 325222 578454
rect 324986 577898 325222 578134
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 324986 506218 325222 506454
rect 324986 505898 325222 506134
rect 324986 470218 325222 470454
rect 324986 469898 325222 470134
rect 317786 427018 318022 427254
rect 317786 426698 318022 426934
rect 317786 391018 318022 391254
rect 317786 390698 318022 390934
rect 317786 355018 318022 355254
rect 317786 354698 318022 354934
rect 317786 319018 318022 319254
rect 317786 318698 318022 318934
rect 317786 283018 318022 283254
rect 317786 282698 318022 282934
rect 317786 247018 318022 247254
rect 317786 246698 318022 246934
rect 317786 211018 318022 211254
rect 317786 210698 318022 210934
rect 317786 175018 318022 175254
rect 317786 174698 318022 174934
rect 317786 139018 318022 139254
rect 317786 138698 318022 138934
rect 317786 103018 318022 103254
rect 317786 102698 318022 102934
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 310586 -3342 310822 -3106
rect 310586 -3662 310822 -3426
rect 314186 -5182 314422 -4946
rect 314186 -5502 314422 -5266
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 324986 398218 325222 398454
rect 324986 397898 325222 398134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 324986 254218 325222 254454
rect 324986 253898 325222 254134
rect 324986 218218 325222 218454
rect 324986 217898 325222 218134
rect 324986 182218 325222 182454
rect 324986 181898 325222 182134
rect 324986 146218 325222 146454
rect 324986 145898 325222 146134
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6102 300022 -5866
rect 299786 -6422 300022 -6186
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 328586 581818 328822 582054
rect 328586 581498 328822 581734
rect 328586 545818 328822 546054
rect 328586 545498 328822 545734
rect 328586 509818 328822 510054
rect 328586 509498 328822 509734
rect 328586 473818 328822 474054
rect 328586 473498 328822 473734
rect 328586 437818 328822 438054
rect 328586 437498 328822 437734
rect 328586 401818 328822 402054
rect 328586 401498 328822 401734
rect 328586 365818 328822 366054
rect 328586 365498 328822 365734
rect 328586 329818 328822 330054
rect 328586 329498 328822 329734
rect 328586 293818 328822 294054
rect 328586 293498 328822 293734
rect 328586 257818 328822 258054
rect 328586 257498 328822 257734
rect 328586 221818 328822 222054
rect 328586 221498 328822 221734
rect 328586 185818 328822 186054
rect 328586 185498 328822 185734
rect 328586 149818 328822 150054
rect 328586 149498 328822 149734
rect 328586 113818 328822 114054
rect 328586 113498 328822 113734
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2422 328822 -2186
rect 328586 -2742 328822 -2506
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 332186 585418 332422 585654
rect 332186 585098 332422 585334
rect 332186 549418 332422 549654
rect 332186 549098 332422 549334
rect 332186 513418 332422 513654
rect 332186 513098 332422 513334
rect 332186 477418 332422 477654
rect 332186 477098 332422 477334
rect 332186 441418 332422 441654
rect 332186 441098 332422 441334
rect 332186 405418 332422 405654
rect 332186 405098 332422 405334
rect 332186 369418 332422 369654
rect 332186 369098 332422 369334
rect 332186 333418 332422 333654
rect 332186 333098 332422 333334
rect 332186 297418 332422 297654
rect 332186 297098 332422 297334
rect 332186 261418 332422 261654
rect 332186 261098 332422 261334
rect 332186 225418 332422 225654
rect 332186 225098 332422 225334
rect 332186 189418 332422 189654
rect 332186 189098 332422 189334
rect 332186 153418 332422 153654
rect 332186 153098 332422 153334
rect 332186 117418 332422 117654
rect 332186 117098 332422 117334
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4262 332422 -4026
rect 332186 -4582 332422 -4346
rect 353786 711042 354022 711278
rect 353786 710722 354022 710958
rect 350186 709202 350422 709438
rect 350186 708882 350422 709118
rect 346586 707362 346822 707598
rect 346586 707042 346822 707278
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 335786 589018 336022 589254
rect 335786 588698 336022 588934
rect 335786 553018 336022 553254
rect 335786 552698 336022 552934
rect 335786 517018 336022 517254
rect 335786 516698 336022 516934
rect 335786 481018 336022 481254
rect 335786 480698 336022 480934
rect 342986 705522 343222 705758
rect 342986 705202 343222 705438
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 342986 560218 343222 560454
rect 342986 559898 343222 560134
rect 342986 524218 343222 524454
rect 342986 523898 343222 524134
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 335786 445018 336022 445254
rect 335786 444698 336022 444934
rect 335786 409018 336022 409254
rect 335786 408698 336022 408934
rect 335786 373018 336022 373254
rect 335786 372698 336022 372934
rect 335786 337018 336022 337254
rect 335786 336698 336022 336934
rect 335786 301018 336022 301254
rect 335786 300698 336022 300934
rect 335786 265018 336022 265254
rect 335786 264698 336022 264934
rect 335786 229018 336022 229254
rect 335786 228698 336022 228934
rect 335786 193018 336022 193254
rect 335786 192698 336022 192934
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 346586 599818 346822 600054
rect 346586 599498 346822 599734
rect 346586 563818 346822 564054
rect 346586 563498 346822 563734
rect 346586 527818 346822 528054
rect 346586 527498 346822 527734
rect 346586 491818 346822 492054
rect 346586 491498 346822 491734
rect 342986 452218 343222 452454
rect 342986 451898 343222 452134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 342986 380218 343222 380454
rect 342986 379898 343222 380134
rect 342986 344218 343222 344454
rect 342986 343898 343222 344134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 342986 272218 343222 272454
rect 342986 271898 343222 272134
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 342986 200218 343222 200454
rect 342986 199898 343222 200134
rect 335786 157018 336022 157254
rect 335786 156698 336022 156934
rect 335786 121018 336022 121254
rect 335786 120698 336022 120934
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 350186 603418 350422 603654
rect 350186 603098 350422 603334
rect 350186 567418 350422 567654
rect 350186 567098 350422 567334
rect 350186 531418 350422 531654
rect 350186 531098 350422 531334
rect 350186 495418 350422 495654
rect 350186 495098 350422 495334
rect 346586 455818 346822 456054
rect 346586 455498 346822 455734
rect 346586 419818 346822 420054
rect 346586 419498 346822 419734
rect 346586 383818 346822 384054
rect 346586 383498 346822 383734
rect 346586 347818 346822 348054
rect 346586 347498 346822 347734
rect 346586 311818 346822 312054
rect 346586 311498 346822 311734
rect 346586 275818 346822 276054
rect 346586 275498 346822 275734
rect 346586 239818 346822 240054
rect 346586 239498 346822 239734
rect 346586 203818 346822 204054
rect 346586 203498 346822 203734
rect 346586 167818 346822 168054
rect 346586 167498 346822 167734
rect 346586 131818 346822 132054
rect 346586 131498 346822 131734
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7022 318022 -6786
rect 317786 -7342 318022 -7106
rect 342986 -1502 343222 -1266
rect 342986 -1822 343222 -1586
rect 350186 459418 350422 459654
rect 350186 459098 350422 459334
rect 350186 423418 350422 423654
rect 350186 423098 350422 423334
rect 350186 387418 350422 387654
rect 350186 387098 350422 387334
rect 350186 351418 350422 351654
rect 350186 351098 350422 351334
rect 350186 315418 350422 315654
rect 350186 315098 350422 315334
rect 350186 279418 350422 279654
rect 350186 279098 350422 279334
rect 350186 243418 350422 243654
rect 350186 243098 350422 243334
rect 350186 207418 350422 207654
rect 350186 207098 350422 207334
rect 350186 171418 350422 171654
rect 350186 171098 350422 171334
rect 350186 135418 350422 135654
rect 350186 135098 350422 135334
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3342 346822 -3106
rect 346586 -3662 346822 -3426
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5182 350422 -4946
rect 350186 -5502 350422 -5266
rect 371786 710122 372022 710358
rect 371786 709802 372022 710038
rect 368186 708282 368422 708518
rect 368186 707962 368422 708198
rect 364586 706442 364822 706678
rect 364586 706122 364822 706358
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 353786 607018 354022 607254
rect 353786 606698 354022 606934
rect 353786 571018 354022 571254
rect 353786 570698 354022 570934
rect 353786 535018 354022 535254
rect 353786 534698 354022 534934
rect 353786 499018 354022 499254
rect 353786 498698 354022 498934
rect 353786 463018 354022 463254
rect 353786 462698 354022 462934
rect 353786 427018 354022 427254
rect 353786 426698 354022 426934
rect 353786 391018 354022 391254
rect 353786 390698 354022 390934
rect 353786 355018 354022 355254
rect 353786 354698 354022 354934
rect 353786 319018 354022 319254
rect 353786 318698 354022 318934
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 360986 578218 361222 578454
rect 360986 577898 361222 578134
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 360986 506218 361222 506454
rect 360986 505898 361222 506134
rect 360986 470218 361222 470454
rect 360986 469898 361222 470134
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 360986 398218 361222 398454
rect 360986 397898 361222 398134
rect 360986 362218 361222 362454
rect 360986 361898 361222 362134
rect 360986 326218 361222 326454
rect 360986 325898 361222 326134
rect 353786 283018 354022 283254
rect 353786 282698 354022 282934
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 353786 247018 354022 247254
rect 353786 246698 354022 246934
rect 360986 254218 361222 254454
rect 360986 253898 361222 254134
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 353786 211018 354022 211254
rect 353786 210698 354022 210934
rect 353786 175018 354022 175254
rect 353786 174698 354022 174934
rect 360986 182218 361222 182454
rect 360986 181898 361222 182134
rect 353786 139018 354022 139254
rect 353786 138698 354022 138934
rect 353786 103018 354022 103254
rect 353786 102698 354022 102934
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6102 336022 -5866
rect 335786 -6422 336022 -6186
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 364586 581818 364822 582054
rect 364586 581498 364822 581734
rect 364586 545818 364822 546054
rect 364586 545498 364822 545734
rect 364586 509818 364822 510054
rect 364586 509498 364822 509734
rect 364586 473818 364822 474054
rect 364586 473498 364822 473734
rect 364586 437818 364822 438054
rect 364586 437498 364822 437734
rect 364586 401818 364822 402054
rect 364586 401498 364822 401734
rect 364586 365818 364822 366054
rect 364586 365498 364822 365734
rect 364586 329818 364822 330054
rect 364586 329498 364822 329734
rect 364586 293818 364822 294054
rect 364586 293498 364822 293734
rect 364586 257818 364822 258054
rect 364586 257498 364822 257734
rect 364586 221818 364822 222054
rect 364586 221498 364822 221734
rect 364586 185818 364822 186054
rect 364586 185498 364822 185734
rect 364586 149818 364822 150054
rect 364586 149498 364822 149734
rect 364586 113818 364822 114054
rect 364586 113498 364822 113734
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 368186 585418 368422 585654
rect 368186 585098 368422 585334
rect 368186 549418 368422 549654
rect 368186 549098 368422 549334
rect 368186 513418 368422 513654
rect 368186 513098 368422 513334
rect 368186 477418 368422 477654
rect 368186 477098 368422 477334
rect 368186 441418 368422 441654
rect 368186 441098 368422 441334
rect 368186 405418 368422 405654
rect 368186 405098 368422 405334
rect 368186 369418 368422 369654
rect 368186 369098 368422 369334
rect 368186 333418 368422 333654
rect 368186 333098 368422 333334
rect 368186 297418 368422 297654
rect 368186 297098 368422 297334
rect 368186 261418 368422 261654
rect 368186 261098 368422 261334
rect 368186 225418 368422 225654
rect 368186 225098 368422 225334
rect 368186 189418 368422 189654
rect 368186 189098 368422 189334
rect 368186 153418 368422 153654
rect 368186 153098 368422 153334
rect 368186 117418 368422 117654
rect 368186 117098 368422 117334
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2422 364822 -2186
rect 364586 -2742 364822 -2506
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4262 368422 -4026
rect 368186 -4582 368422 -4346
rect 389786 711042 390022 711278
rect 389786 710722 390022 710958
rect 386186 709202 386422 709438
rect 386186 708882 386422 709118
rect 382586 707362 382822 707598
rect 382586 707042 382822 707278
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 371786 589018 372022 589254
rect 371786 588698 372022 588934
rect 371786 553018 372022 553254
rect 371786 552698 372022 552934
rect 371786 517018 372022 517254
rect 371786 516698 372022 516934
rect 371786 481018 372022 481254
rect 371786 480698 372022 480934
rect 371786 445018 372022 445254
rect 371786 444698 372022 444934
rect 371786 409018 372022 409254
rect 371786 408698 372022 408934
rect 371786 373018 372022 373254
rect 371786 372698 372022 372934
rect 371786 337018 372022 337254
rect 371786 336698 372022 336934
rect 378986 705522 379222 705758
rect 378986 705202 379222 705438
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 378986 452218 379222 452454
rect 378986 451898 379222 452134
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 378986 380218 379222 380454
rect 378986 379898 379222 380134
rect 378986 344218 379222 344454
rect 378986 343898 379222 344134
rect 371786 301018 372022 301254
rect 371786 300698 372022 300934
rect 371786 265018 372022 265254
rect 371786 264698 372022 264934
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 378986 272218 379222 272454
rect 378986 271898 379222 272134
rect 371786 229018 372022 229254
rect 371786 228698 372022 228934
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 371786 193018 372022 193254
rect 371786 192698 372022 192934
rect 378986 200218 379222 200454
rect 378986 199898 379222 200134
rect 371786 157018 372022 157254
rect 371786 156698 372022 156934
rect 371786 121018 372022 121254
rect 371786 120698 372022 120934
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7022 354022 -6786
rect 353786 -7342 354022 -7106
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1502 379222 -1266
rect 378986 -1822 379222 -1586
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 382586 599818 382822 600054
rect 382586 599498 382822 599734
rect 382586 563818 382822 564054
rect 382586 563498 382822 563734
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 382586 491818 382822 492054
rect 382586 491498 382822 491734
rect 382586 455818 382822 456054
rect 382586 455498 382822 455734
rect 382586 419818 382822 420054
rect 382586 419498 382822 419734
rect 382586 383818 382822 384054
rect 382586 383498 382822 383734
rect 382586 347818 382822 348054
rect 382586 347498 382822 347734
rect 382586 311818 382822 312054
rect 382586 311498 382822 311734
rect 382586 275818 382822 276054
rect 382586 275498 382822 275734
rect 382586 239818 382822 240054
rect 382586 239498 382822 239734
rect 382586 203818 382822 204054
rect 382586 203498 382822 203734
rect 382586 167818 382822 168054
rect 382586 167498 382822 167734
rect 382586 131818 382822 132054
rect 382586 131498 382822 131734
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3342 382822 -3106
rect 382586 -3662 382822 -3426
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 386186 639418 386422 639654
rect 386186 639098 386422 639334
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 386186 567418 386422 567654
rect 386186 567098 386422 567334
rect 386186 531418 386422 531654
rect 386186 531098 386422 531334
rect 386186 495418 386422 495654
rect 386186 495098 386422 495334
rect 386186 459418 386422 459654
rect 386186 459098 386422 459334
rect 386186 423418 386422 423654
rect 386186 423098 386422 423334
rect 386186 387418 386422 387654
rect 386186 387098 386422 387334
rect 386186 351418 386422 351654
rect 386186 351098 386422 351334
rect 386186 315418 386422 315654
rect 386186 315098 386422 315334
rect 386186 279418 386422 279654
rect 386186 279098 386422 279334
rect 386186 243418 386422 243654
rect 386186 243098 386422 243334
rect 386186 207418 386422 207654
rect 386186 207098 386422 207334
rect 386186 171418 386422 171654
rect 386186 171098 386422 171334
rect 386186 135418 386422 135654
rect 386186 135098 386422 135334
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5182 386422 -4946
rect 386186 -5502 386422 -5266
rect 407786 710122 408022 710358
rect 407786 709802 408022 710038
rect 404186 708282 404422 708518
rect 404186 707962 404422 708198
rect 400586 706442 400822 706678
rect 400586 706122 400822 706358
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 389786 571018 390022 571254
rect 389786 570698 390022 570934
rect 389786 535018 390022 535254
rect 389786 534698 390022 534934
rect 389786 499018 390022 499254
rect 389786 498698 390022 498934
rect 389786 463018 390022 463254
rect 389786 462698 390022 462934
rect 389786 427018 390022 427254
rect 389786 426698 390022 426934
rect 389786 391018 390022 391254
rect 389786 390698 390022 390934
rect 389786 355018 390022 355254
rect 389786 354698 390022 354934
rect 389786 319018 390022 319254
rect 389786 318698 390022 318934
rect 389786 283018 390022 283254
rect 389786 282698 390022 282934
rect 389786 247018 390022 247254
rect 389786 246698 390022 246934
rect 389786 211018 390022 211254
rect 389786 210698 390022 210934
rect 389786 175018 390022 175254
rect 389786 174698 390022 174934
rect 389786 139018 390022 139254
rect 389786 138698 390022 138934
rect 389786 103018 390022 103254
rect 389786 102698 390022 102934
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6102 372022 -5866
rect 371786 -6422 372022 -6186
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 396986 470218 397222 470454
rect 396986 469898 397222 470134
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 396986 398218 397222 398454
rect 396986 397898 397222 398134
rect 396986 362218 397222 362454
rect 396986 361898 397222 362134
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 396986 254218 397222 254454
rect 396986 253898 397222 254134
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 400586 509818 400822 510054
rect 400586 509498 400822 509734
rect 400586 473818 400822 474054
rect 400586 473498 400822 473734
rect 400586 437818 400822 438054
rect 400586 437498 400822 437734
rect 400586 401818 400822 402054
rect 400586 401498 400822 401734
rect 400586 365818 400822 366054
rect 400586 365498 400822 365734
rect 400586 329818 400822 330054
rect 400586 329498 400822 329734
rect 400586 293818 400822 294054
rect 400586 293498 400822 293734
rect 400586 257818 400822 258054
rect 400586 257498 400822 257734
rect 400586 221818 400822 222054
rect 400586 221498 400822 221734
rect 400586 185818 400822 186054
rect 400586 185498 400822 185734
rect 400586 149818 400822 150054
rect 400586 149498 400822 149734
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2422 400822 -2186
rect 400586 -2742 400822 -2506
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 404186 513418 404422 513654
rect 404186 513098 404422 513334
rect 404186 477418 404422 477654
rect 404186 477098 404422 477334
rect 404186 441418 404422 441654
rect 404186 441098 404422 441334
rect 404186 405418 404422 405654
rect 404186 405098 404422 405334
rect 404186 369418 404422 369654
rect 404186 369098 404422 369334
rect 404186 333418 404422 333654
rect 404186 333098 404422 333334
rect 404186 297418 404422 297654
rect 404186 297098 404422 297334
rect 404186 261418 404422 261654
rect 404186 261098 404422 261334
rect 404186 225418 404422 225654
rect 404186 225098 404422 225334
rect 404186 189418 404422 189654
rect 404186 189098 404422 189334
rect 404186 153418 404422 153654
rect 404186 153098 404422 153334
rect 404186 117418 404422 117654
rect 404186 117098 404422 117334
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4262 404422 -4026
rect 404186 -4582 404422 -4346
rect 425786 711042 426022 711278
rect 425786 710722 426022 710958
rect 422186 709202 422422 709438
rect 422186 708882 422422 709118
rect 418586 707362 418822 707598
rect 418586 707042 418822 707278
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 407786 517018 408022 517254
rect 407786 516698 408022 516934
rect 407786 481018 408022 481254
rect 407786 480698 408022 480934
rect 407786 445018 408022 445254
rect 407786 444698 408022 444934
rect 407786 409018 408022 409254
rect 407786 408698 408022 408934
rect 407786 373018 408022 373254
rect 407786 372698 408022 372934
rect 407786 337018 408022 337254
rect 407786 336698 408022 336934
rect 407786 301018 408022 301254
rect 407786 300698 408022 300934
rect 407786 265018 408022 265254
rect 407786 264698 408022 264934
rect 407786 229018 408022 229254
rect 407786 228698 408022 228934
rect 407786 193018 408022 193254
rect 407786 192698 408022 192934
rect 407786 157018 408022 157254
rect 407786 156698 408022 156934
rect 407786 121018 408022 121254
rect 407786 120698 408022 120934
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7022 390022 -6786
rect 389786 -7342 390022 -7106
rect 414986 705522 415222 705758
rect 414986 705202 415222 705438
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1502 415222 -1266
rect 414986 -1822 415222 -1586
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 418586 527818 418822 528054
rect 418586 527498 418822 527734
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 418586 455818 418822 456054
rect 418586 455498 418822 455734
rect 418586 419818 418822 420054
rect 418586 419498 418822 419734
rect 418586 383818 418822 384054
rect 418586 383498 418822 383734
rect 418586 347818 418822 348054
rect 418586 347498 418822 347734
rect 418586 311818 418822 312054
rect 418586 311498 418822 311734
rect 418586 275818 418822 276054
rect 418586 275498 418822 275734
rect 418586 239818 418822 240054
rect 418586 239498 418822 239734
rect 418586 203818 418822 204054
rect 418586 203498 418822 203734
rect 418586 167818 418822 168054
rect 418586 167498 418822 167734
rect 418586 131818 418822 132054
rect 418586 131498 418822 131734
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3342 418822 -3106
rect 418586 -3662 418822 -3426
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 422186 567418 422422 567654
rect 422186 567098 422422 567334
rect 422186 531418 422422 531654
rect 422186 531098 422422 531334
rect 422186 495418 422422 495654
rect 422186 495098 422422 495334
rect 422186 459418 422422 459654
rect 422186 459098 422422 459334
rect 422186 423418 422422 423654
rect 422186 423098 422422 423334
rect 422186 387418 422422 387654
rect 422186 387098 422422 387334
rect 422186 351418 422422 351654
rect 422186 351098 422422 351334
rect 422186 315418 422422 315654
rect 422186 315098 422422 315334
rect 422186 279418 422422 279654
rect 422186 279098 422422 279334
rect 422186 243418 422422 243654
rect 422186 243098 422422 243334
rect 422186 207418 422422 207654
rect 422186 207098 422422 207334
rect 422186 171418 422422 171654
rect 422186 171098 422422 171334
rect 422186 135418 422422 135654
rect 422186 135098 422422 135334
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5182 422422 -4946
rect 422186 -5502 422422 -5266
rect 443786 710122 444022 710358
rect 443786 709802 444022 710038
rect 440186 708282 440422 708518
rect 440186 707962 440422 708198
rect 436586 706442 436822 706678
rect 436586 706122 436822 706358
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 425786 571018 426022 571254
rect 425786 570698 426022 570934
rect 425786 535018 426022 535254
rect 425786 534698 426022 534934
rect 425786 499018 426022 499254
rect 425786 498698 426022 498934
rect 425786 463018 426022 463254
rect 425786 462698 426022 462934
rect 425786 427018 426022 427254
rect 425786 426698 426022 426934
rect 425786 391018 426022 391254
rect 425786 390698 426022 390934
rect 425786 355018 426022 355254
rect 425786 354698 426022 354934
rect 425786 319018 426022 319254
rect 425786 318698 426022 318934
rect 425786 283018 426022 283254
rect 425786 282698 426022 282934
rect 425786 247018 426022 247254
rect 425786 246698 426022 246934
rect 425786 211018 426022 211254
rect 425786 210698 426022 210934
rect 425786 175018 426022 175254
rect 425786 174698 426022 174934
rect 425786 139018 426022 139254
rect 425786 138698 426022 138934
rect 425786 103018 426022 103254
rect 425786 102698 426022 102934
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6102 408022 -5866
rect 407786 -6422 408022 -6186
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 436586 581818 436822 582054
rect 436586 581498 436822 581734
rect 436586 545818 436822 546054
rect 436586 545498 436822 545734
rect 436586 509818 436822 510054
rect 436586 509498 436822 509734
rect 436586 473818 436822 474054
rect 436586 473498 436822 473734
rect 436586 437818 436822 438054
rect 436586 437498 436822 437734
rect 436586 401818 436822 402054
rect 436586 401498 436822 401734
rect 436586 365818 436822 366054
rect 436586 365498 436822 365734
rect 436586 329818 436822 330054
rect 436586 329498 436822 329734
rect 436586 293818 436822 294054
rect 436586 293498 436822 293734
rect 436586 257818 436822 258054
rect 436586 257498 436822 257734
rect 436586 221818 436822 222054
rect 436586 221498 436822 221734
rect 436586 185818 436822 186054
rect 436586 185498 436822 185734
rect 436586 149818 436822 150054
rect 436586 149498 436822 149734
rect 436586 113818 436822 114054
rect 436586 113498 436822 113734
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2422 436822 -2186
rect 436586 -2742 436822 -2506
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 440186 585418 440422 585654
rect 440186 585098 440422 585334
rect 440186 549418 440422 549654
rect 440186 549098 440422 549334
rect 440186 513418 440422 513654
rect 440186 513098 440422 513334
rect 440186 477418 440422 477654
rect 440186 477098 440422 477334
rect 440186 441418 440422 441654
rect 440186 441098 440422 441334
rect 440186 405418 440422 405654
rect 440186 405098 440422 405334
rect 440186 369418 440422 369654
rect 440186 369098 440422 369334
rect 440186 333418 440422 333654
rect 440186 333098 440422 333334
rect 440186 297418 440422 297654
rect 440186 297098 440422 297334
rect 440186 261418 440422 261654
rect 440186 261098 440422 261334
rect 440186 225418 440422 225654
rect 440186 225098 440422 225334
rect 440186 189418 440422 189654
rect 440186 189098 440422 189334
rect 440186 153418 440422 153654
rect 440186 153098 440422 153334
rect 440186 117418 440422 117654
rect 440186 117098 440422 117334
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4262 440422 -4026
rect 440186 -4582 440422 -4346
rect 461786 711042 462022 711278
rect 461786 710722 462022 710958
rect 458186 709202 458422 709438
rect 458186 708882 458422 709118
rect 454586 707362 454822 707598
rect 454586 707042 454822 707278
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 443786 589018 444022 589254
rect 443786 588698 444022 588934
rect 443786 553018 444022 553254
rect 443786 552698 444022 552934
rect 443786 517018 444022 517254
rect 443786 516698 444022 516934
rect 443786 481018 444022 481254
rect 443786 480698 444022 480934
rect 443786 445018 444022 445254
rect 443786 444698 444022 444934
rect 443786 409018 444022 409254
rect 443786 408698 444022 408934
rect 443786 373018 444022 373254
rect 443786 372698 444022 372934
rect 443786 337018 444022 337254
rect 443786 336698 444022 336934
rect 443786 301018 444022 301254
rect 443786 300698 444022 300934
rect 443786 265018 444022 265254
rect 443786 264698 444022 264934
rect 443786 229018 444022 229254
rect 443786 228698 444022 228934
rect 443786 193018 444022 193254
rect 443786 192698 444022 192934
rect 443786 157018 444022 157254
rect 443786 156698 444022 156934
rect 443786 121018 444022 121254
rect 443786 120698 444022 120934
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7022 426022 -6786
rect 425786 -7342 426022 -7106
rect 450986 705522 451222 705758
rect 450986 705202 451222 705438
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1502 451222 -1266
rect 450986 -1822 451222 -1586
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 454586 599818 454822 600054
rect 454586 599498 454822 599734
rect 454586 563818 454822 564054
rect 454586 563498 454822 563734
rect 454586 527818 454822 528054
rect 454586 527498 454822 527734
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 454586 383818 454822 384054
rect 454586 383498 454822 383734
rect 454586 347818 454822 348054
rect 454586 347498 454822 347734
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 454586 275818 454822 276054
rect 454586 275498 454822 275734
rect 454586 239818 454822 240054
rect 454586 239498 454822 239734
rect 454586 203818 454822 204054
rect 454586 203498 454822 203734
rect 454586 167818 454822 168054
rect 454586 167498 454822 167734
rect 454586 131818 454822 132054
rect 454586 131498 454822 131734
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3342 454822 -3106
rect 454586 -3662 454822 -3426
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 458186 603418 458422 603654
rect 458186 603098 458422 603334
rect 458186 567418 458422 567654
rect 458186 567098 458422 567334
rect 458186 531418 458422 531654
rect 458186 531098 458422 531334
rect 458186 495418 458422 495654
rect 458186 495098 458422 495334
rect 458186 459418 458422 459654
rect 458186 459098 458422 459334
rect 458186 423418 458422 423654
rect 458186 423098 458422 423334
rect 458186 387418 458422 387654
rect 458186 387098 458422 387334
rect 458186 351418 458422 351654
rect 458186 351098 458422 351334
rect 458186 315418 458422 315654
rect 458186 315098 458422 315334
rect 458186 279418 458422 279654
rect 458186 279098 458422 279334
rect 458186 243418 458422 243654
rect 458186 243098 458422 243334
rect 458186 207418 458422 207654
rect 458186 207098 458422 207334
rect 458186 171418 458422 171654
rect 458186 171098 458422 171334
rect 458186 135418 458422 135654
rect 458186 135098 458422 135334
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5182 458422 -4946
rect 458186 -5502 458422 -5266
rect 479786 710122 480022 710358
rect 479786 709802 480022 710038
rect 476186 708282 476422 708518
rect 476186 707962 476422 708198
rect 472586 706442 472822 706678
rect 472586 706122 472822 706358
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 461786 607018 462022 607254
rect 461786 606698 462022 606934
rect 461786 571018 462022 571254
rect 461786 570698 462022 570934
rect 461786 535018 462022 535254
rect 461786 534698 462022 534934
rect 461786 499018 462022 499254
rect 461786 498698 462022 498934
rect 461786 463018 462022 463254
rect 461786 462698 462022 462934
rect 461786 427018 462022 427254
rect 461786 426698 462022 426934
rect 461786 391018 462022 391254
rect 461786 390698 462022 390934
rect 461786 355018 462022 355254
rect 461786 354698 462022 354934
rect 461786 319018 462022 319254
rect 461786 318698 462022 318934
rect 461786 283018 462022 283254
rect 461786 282698 462022 282934
rect 461786 247018 462022 247254
rect 461786 246698 462022 246934
rect 461786 211018 462022 211254
rect 461786 210698 462022 210934
rect 461786 175018 462022 175254
rect 461786 174698 462022 174934
rect 461786 139018 462022 139254
rect 461786 138698 462022 138934
rect 461786 103018 462022 103254
rect 461786 102698 462022 102934
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6102 444022 -5866
rect 443786 -6422 444022 -6186
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 472586 581818 472822 582054
rect 472586 581498 472822 581734
rect 472586 545818 472822 546054
rect 472586 545498 472822 545734
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 472586 473818 472822 474054
rect 472586 473498 472822 473734
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 472586 401818 472822 402054
rect 472586 401498 472822 401734
rect 472586 365818 472822 366054
rect 472586 365498 472822 365734
rect 472586 329818 472822 330054
rect 472586 329498 472822 329734
rect 472586 293818 472822 294054
rect 472586 293498 472822 293734
rect 472586 257818 472822 258054
rect 472586 257498 472822 257734
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 472586 185818 472822 186054
rect 472586 185498 472822 185734
rect 472586 149818 472822 150054
rect 472586 149498 472822 149734
rect 472586 113818 472822 114054
rect 472586 113498 472822 113734
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2422 472822 -2186
rect 472586 -2742 472822 -2506
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 476186 585418 476422 585654
rect 476186 585098 476422 585334
rect 476186 549418 476422 549654
rect 476186 549098 476422 549334
rect 476186 513418 476422 513654
rect 476186 513098 476422 513334
rect 476186 477418 476422 477654
rect 476186 477098 476422 477334
rect 476186 441418 476422 441654
rect 476186 441098 476422 441334
rect 476186 405418 476422 405654
rect 476186 405098 476422 405334
rect 476186 369418 476422 369654
rect 476186 369098 476422 369334
rect 476186 333418 476422 333654
rect 476186 333098 476422 333334
rect 476186 297418 476422 297654
rect 476186 297098 476422 297334
rect 476186 261418 476422 261654
rect 476186 261098 476422 261334
rect 476186 225418 476422 225654
rect 476186 225098 476422 225334
rect 476186 189418 476422 189654
rect 476186 189098 476422 189334
rect 476186 153418 476422 153654
rect 476186 153098 476422 153334
rect 476186 117418 476422 117654
rect 476186 117098 476422 117334
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4262 476422 -4026
rect 476186 -4582 476422 -4346
rect 497786 711042 498022 711278
rect 497786 710722 498022 710958
rect 494186 709202 494422 709438
rect 494186 708882 494422 709118
rect 490586 707362 490822 707598
rect 490586 707042 490822 707278
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 479786 589018 480022 589254
rect 479786 588698 480022 588934
rect 479786 553018 480022 553254
rect 479786 552698 480022 552934
rect 479786 517018 480022 517254
rect 479786 516698 480022 516934
rect 479786 481018 480022 481254
rect 479786 480698 480022 480934
rect 479786 445018 480022 445254
rect 479786 444698 480022 444934
rect 479786 409018 480022 409254
rect 479786 408698 480022 408934
rect 479786 373018 480022 373254
rect 479786 372698 480022 372934
rect 479786 337018 480022 337254
rect 479786 336698 480022 336934
rect 479786 301018 480022 301254
rect 479786 300698 480022 300934
rect 479786 265018 480022 265254
rect 479786 264698 480022 264934
rect 479786 229018 480022 229254
rect 479786 228698 480022 228934
rect 479786 193018 480022 193254
rect 479786 192698 480022 192934
rect 479786 157018 480022 157254
rect 479786 156698 480022 156934
rect 479786 121018 480022 121254
rect 479786 120698 480022 120934
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 486986 705522 487222 705758
rect 486986 705202 487222 705438
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7022 462022 -6786
rect 461786 -7342 462022 -7106
rect 486986 -1502 487222 -1266
rect 486986 -1822 487222 -1586
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 490586 599818 490822 600054
rect 490586 599498 490822 599734
rect 490586 563818 490822 564054
rect 490586 563498 490822 563734
rect 490586 527818 490822 528054
rect 490586 527498 490822 527734
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 490586 383818 490822 384054
rect 490586 383498 490822 383734
rect 490586 347818 490822 348054
rect 490586 347498 490822 347734
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 490586 275818 490822 276054
rect 490586 275498 490822 275734
rect 490586 239818 490822 240054
rect 490586 239498 490822 239734
rect 490586 203818 490822 204054
rect 490586 203498 490822 203734
rect 490586 167818 490822 168054
rect 490586 167498 490822 167734
rect 490586 131818 490822 132054
rect 490586 131498 490822 131734
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3342 490822 -3106
rect 490586 -3662 490822 -3426
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 494186 603418 494422 603654
rect 494186 603098 494422 603334
rect 494186 567418 494422 567654
rect 494186 567098 494422 567334
rect 494186 531418 494422 531654
rect 494186 531098 494422 531334
rect 494186 495418 494422 495654
rect 494186 495098 494422 495334
rect 494186 459418 494422 459654
rect 494186 459098 494422 459334
rect 494186 423418 494422 423654
rect 494186 423098 494422 423334
rect 494186 387418 494422 387654
rect 494186 387098 494422 387334
rect 494186 351418 494422 351654
rect 494186 351098 494422 351334
rect 494186 315418 494422 315654
rect 494186 315098 494422 315334
rect 494186 279418 494422 279654
rect 494186 279098 494422 279334
rect 494186 243418 494422 243654
rect 494186 243098 494422 243334
rect 494186 207418 494422 207654
rect 494186 207098 494422 207334
rect 494186 171418 494422 171654
rect 494186 171098 494422 171334
rect 494186 135418 494422 135654
rect 494186 135098 494422 135334
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5182 494422 -4946
rect 494186 -5502 494422 -5266
rect 515786 710122 516022 710358
rect 515786 709802 516022 710038
rect 512186 708282 512422 708518
rect 512186 707962 512422 708198
rect 508586 706442 508822 706678
rect 508586 706122 508822 706358
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 497786 607018 498022 607254
rect 497786 606698 498022 606934
rect 497786 571018 498022 571254
rect 497786 570698 498022 570934
rect 497786 535018 498022 535254
rect 497786 534698 498022 534934
rect 497786 499018 498022 499254
rect 497786 498698 498022 498934
rect 497786 463018 498022 463254
rect 497786 462698 498022 462934
rect 497786 427018 498022 427254
rect 497786 426698 498022 426934
rect 497786 391018 498022 391254
rect 497786 390698 498022 390934
rect 497786 355018 498022 355254
rect 497786 354698 498022 354934
rect 497786 319018 498022 319254
rect 497786 318698 498022 318934
rect 497786 283018 498022 283254
rect 497786 282698 498022 282934
rect 497786 247018 498022 247254
rect 497786 246698 498022 246934
rect 497786 211018 498022 211254
rect 497786 210698 498022 210934
rect 497786 175018 498022 175254
rect 497786 174698 498022 174934
rect 497786 139018 498022 139254
rect 497786 138698 498022 138934
rect 497786 103018 498022 103254
rect 497786 102698 498022 102934
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6102 480022 -5866
rect 479786 -6422 480022 -6186
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2422 508822 -2186
rect 508586 -2742 508822 -2506
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4262 512422 -4026
rect 512186 -4582 512422 -4346
rect 533786 711042 534022 711278
rect 533786 710722 534022 710958
rect 530186 709202 530422 709438
rect 530186 708882 530422 709118
rect 526586 707362 526822 707598
rect 526586 707042 526822 707278
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7022 498022 -6786
rect 497786 -7342 498022 -7106
rect 522986 705522 523222 705758
rect 522986 705202 523222 705438
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1502 523222 -1266
rect 522986 -1822 523222 -1586
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3342 526822 -3106
rect 526586 -3662 526822 -3426
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5182 530422 -4946
rect 530186 -5502 530422 -5266
rect 551786 710122 552022 710358
rect 551786 709802 552022 710038
rect 548186 708282 548422 708518
rect 548186 707962 548422 708198
rect 544586 706442 544822 706678
rect 544586 706122 544822 706358
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6102 516022 -5866
rect 515786 -6422 516022 -6186
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2422 544822 -2186
rect 544586 -2742 544822 -2506
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4262 548422 -4026
rect 548186 -4582 548422 -4346
rect 569786 711042 570022 711278
rect 569786 710722 570022 710958
rect 566186 709202 566422 709438
rect 566186 708882 566422 709118
rect 562586 707362 562822 707598
rect 562586 707042 562822 707278
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7022 534022 -6786
rect 533786 -7342 534022 -7106
rect 558986 705522 559222 705758
rect 558986 705202 559222 705438
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1502 559222 -1266
rect 558986 -1822 559222 -1586
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3342 562822 -3106
rect 562586 -3662 562822 -3426
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5182 566422 -4946
rect 566186 -5502 566422 -5266
rect 591942 711042 592178 711278
rect 591942 710722 592178 710958
rect 591022 710122 591258 710358
rect 591022 709802 591258 710038
rect 590102 709202 590338 709438
rect 590102 708882 590338 709118
rect 589182 708282 589418 708518
rect 589182 707962 589418 708198
rect 588262 707362 588498 707598
rect 588262 707042 588498 707278
rect 580586 706442 580822 706678
rect 580586 706122 580822 706358
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6102 552022 -5866
rect 551786 -6422 552022 -6186
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587342 706442 587578 706678
rect 587342 706122 587578 706358
rect 586422 705522 586658 705758
rect 586422 705202 586658 705438
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586422 668218 586658 668454
rect 586422 667898 586658 668134
rect 586422 632218 586658 632454
rect 586422 631898 586658 632134
rect 586422 596218 586658 596454
rect 586422 595898 586658 596134
rect 586422 560218 586658 560454
rect 586422 559898 586658 560134
rect 586422 524218 586658 524454
rect 586422 523898 586658 524134
rect 586422 488218 586658 488454
rect 586422 487898 586658 488134
rect 586422 452218 586658 452454
rect 586422 451898 586658 452134
rect 586422 416218 586658 416454
rect 586422 415898 586658 416134
rect 586422 380218 586658 380454
rect 586422 379898 586658 380134
rect 586422 344218 586658 344454
rect 586422 343898 586658 344134
rect 586422 308218 586658 308454
rect 586422 307898 586658 308134
rect 586422 272218 586658 272454
rect 586422 271898 586658 272134
rect 586422 236218 586658 236454
rect 586422 235898 586658 236134
rect 586422 200218 586658 200454
rect 586422 199898 586658 200134
rect 586422 164218 586658 164454
rect 586422 163898 586658 164134
rect 586422 128218 586658 128454
rect 586422 127898 586658 128134
rect 586422 92218 586658 92454
rect 586422 91898 586658 92134
rect 586422 56218 586658 56454
rect 586422 55898 586658 56134
rect 586422 20218 586658 20454
rect 586422 19898 586658 20134
rect 586422 -1502 586658 -1266
rect 586422 -1822 586658 -1586
rect 587342 689818 587578 690054
rect 587342 689498 587578 689734
rect 587342 653818 587578 654054
rect 587342 653498 587578 653734
rect 587342 617818 587578 618054
rect 587342 617498 587578 617734
rect 587342 581818 587578 582054
rect 587342 581498 587578 581734
rect 587342 545818 587578 546054
rect 587342 545498 587578 545734
rect 587342 509818 587578 510054
rect 587342 509498 587578 509734
rect 587342 473818 587578 474054
rect 587342 473498 587578 473734
rect 587342 437818 587578 438054
rect 587342 437498 587578 437734
rect 587342 401818 587578 402054
rect 587342 401498 587578 401734
rect 587342 365818 587578 366054
rect 587342 365498 587578 365734
rect 587342 329818 587578 330054
rect 587342 329498 587578 329734
rect 587342 293818 587578 294054
rect 587342 293498 587578 293734
rect 587342 257818 587578 258054
rect 587342 257498 587578 257734
rect 587342 221818 587578 222054
rect 587342 221498 587578 221734
rect 587342 185818 587578 186054
rect 587342 185498 587578 185734
rect 587342 149818 587578 150054
rect 587342 149498 587578 149734
rect 587342 113818 587578 114054
rect 587342 113498 587578 113734
rect 587342 77818 587578 78054
rect 587342 77498 587578 77734
rect 587342 41818 587578 42054
rect 587342 41498 587578 41734
rect 587342 5818 587578 6054
rect 587342 5498 587578 5734
rect 580586 -2422 580822 -2186
rect 580586 -2742 580822 -2506
rect 587342 -2422 587578 -2186
rect 587342 -2742 587578 -2506
rect 588262 671818 588498 672054
rect 588262 671498 588498 671734
rect 588262 635818 588498 636054
rect 588262 635498 588498 635734
rect 588262 599818 588498 600054
rect 588262 599498 588498 599734
rect 588262 563818 588498 564054
rect 588262 563498 588498 563734
rect 588262 527818 588498 528054
rect 588262 527498 588498 527734
rect 588262 491818 588498 492054
rect 588262 491498 588498 491734
rect 588262 455818 588498 456054
rect 588262 455498 588498 455734
rect 588262 419818 588498 420054
rect 588262 419498 588498 419734
rect 588262 383818 588498 384054
rect 588262 383498 588498 383734
rect 588262 347818 588498 348054
rect 588262 347498 588498 347734
rect 588262 311818 588498 312054
rect 588262 311498 588498 311734
rect 588262 275818 588498 276054
rect 588262 275498 588498 275734
rect 588262 239818 588498 240054
rect 588262 239498 588498 239734
rect 588262 203818 588498 204054
rect 588262 203498 588498 203734
rect 588262 167818 588498 168054
rect 588262 167498 588498 167734
rect 588262 131818 588498 132054
rect 588262 131498 588498 131734
rect 588262 95818 588498 96054
rect 588262 95498 588498 95734
rect 588262 59818 588498 60054
rect 588262 59498 588498 59734
rect 588262 23818 588498 24054
rect 588262 23498 588498 23734
rect 588262 -3342 588498 -3106
rect 588262 -3662 588498 -3426
rect 589182 693418 589418 693654
rect 589182 693098 589418 693334
rect 589182 657418 589418 657654
rect 589182 657098 589418 657334
rect 589182 621418 589418 621654
rect 589182 621098 589418 621334
rect 589182 585418 589418 585654
rect 589182 585098 589418 585334
rect 589182 549418 589418 549654
rect 589182 549098 589418 549334
rect 589182 513418 589418 513654
rect 589182 513098 589418 513334
rect 589182 477418 589418 477654
rect 589182 477098 589418 477334
rect 589182 441418 589418 441654
rect 589182 441098 589418 441334
rect 589182 405418 589418 405654
rect 589182 405098 589418 405334
rect 589182 369418 589418 369654
rect 589182 369098 589418 369334
rect 589182 333418 589418 333654
rect 589182 333098 589418 333334
rect 589182 297418 589418 297654
rect 589182 297098 589418 297334
rect 589182 261418 589418 261654
rect 589182 261098 589418 261334
rect 589182 225418 589418 225654
rect 589182 225098 589418 225334
rect 589182 189418 589418 189654
rect 589182 189098 589418 189334
rect 589182 153418 589418 153654
rect 589182 153098 589418 153334
rect 589182 117418 589418 117654
rect 589182 117098 589418 117334
rect 589182 81418 589418 81654
rect 589182 81098 589418 81334
rect 589182 45418 589418 45654
rect 589182 45098 589418 45334
rect 589182 9418 589418 9654
rect 589182 9098 589418 9334
rect 589182 -4262 589418 -4026
rect 589182 -4582 589418 -4346
rect 590102 675418 590338 675654
rect 590102 675098 590338 675334
rect 590102 639418 590338 639654
rect 590102 639098 590338 639334
rect 590102 603418 590338 603654
rect 590102 603098 590338 603334
rect 590102 567418 590338 567654
rect 590102 567098 590338 567334
rect 590102 531418 590338 531654
rect 590102 531098 590338 531334
rect 590102 495418 590338 495654
rect 590102 495098 590338 495334
rect 590102 459418 590338 459654
rect 590102 459098 590338 459334
rect 590102 423418 590338 423654
rect 590102 423098 590338 423334
rect 590102 387418 590338 387654
rect 590102 387098 590338 387334
rect 590102 351418 590338 351654
rect 590102 351098 590338 351334
rect 590102 315418 590338 315654
rect 590102 315098 590338 315334
rect 590102 279418 590338 279654
rect 590102 279098 590338 279334
rect 590102 243418 590338 243654
rect 590102 243098 590338 243334
rect 590102 207418 590338 207654
rect 590102 207098 590338 207334
rect 590102 171418 590338 171654
rect 590102 171098 590338 171334
rect 590102 135418 590338 135654
rect 590102 135098 590338 135334
rect 590102 99418 590338 99654
rect 590102 99098 590338 99334
rect 590102 63418 590338 63654
rect 590102 63098 590338 63334
rect 590102 27418 590338 27654
rect 590102 27098 590338 27334
rect 590102 -5182 590338 -4946
rect 590102 -5502 590338 -5266
rect 591022 697018 591258 697254
rect 591022 696698 591258 696934
rect 591022 661018 591258 661254
rect 591022 660698 591258 660934
rect 591022 625018 591258 625254
rect 591022 624698 591258 624934
rect 591022 589018 591258 589254
rect 591022 588698 591258 588934
rect 591022 553018 591258 553254
rect 591022 552698 591258 552934
rect 591022 517018 591258 517254
rect 591022 516698 591258 516934
rect 591022 481018 591258 481254
rect 591022 480698 591258 480934
rect 591022 445018 591258 445254
rect 591022 444698 591258 444934
rect 591022 409018 591258 409254
rect 591022 408698 591258 408934
rect 591022 373018 591258 373254
rect 591022 372698 591258 372934
rect 591022 337018 591258 337254
rect 591022 336698 591258 336934
rect 591022 301018 591258 301254
rect 591022 300698 591258 300934
rect 591022 265018 591258 265254
rect 591022 264698 591258 264934
rect 591022 229018 591258 229254
rect 591022 228698 591258 228934
rect 591022 193018 591258 193254
rect 591022 192698 591258 192934
rect 591022 157018 591258 157254
rect 591022 156698 591258 156934
rect 591022 121018 591258 121254
rect 591022 120698 591258 120934
rect 591022 85018 591258 85254
rect 591022 84698 591258 84934
rect 591022 49018 591258 49254
rect 591022 48698 591258 48934
rect 591022 13018 591258 13254
rect 591022 12698 591258 12934
rect 591022 -6102 591258 -5866
rect 591022 -6422 591258 -6186
rect 591942 679018 592178 679254
rect 591942 678698 592178 678934
rect 591942 643018 592178 643254
rect 591942 642698 592178 642934
rect 591942 607018 592178 607254
rect 591942 606698 592178 606934
rect 591942 571018 592178 571254
rect 591942 570698 592178 570934
rect 591942 535018 592178 535254
rect 591942 534698 592178 534934
rect 591942 499018 592178 499254
rect 591942 498698 592178 498934
rect 591942 463018 592178 463254
rect 591942 462698 592178 462934
rect 591942 427018 592178 427254
rect 591942 426698 592178 426934
rect 591942 391018 592178 391254
rect 591942 390698 592178 390934
rect 591942 355018 592178 355254
rect 591942 354698 592178 354934
rect 591942 319018 592178 319254
rect 591942 318698 592178 318934
rect 591942 283018 592178 283254
rect 591942 282698 592178 282934
rect 591942 247018 592178 247254
rect 591942 246698 592178 246934
rect 591942 211018 592178 211254
rect 591942 210698 592178 210934
rect 591942 175018 592178 175254
rect 591942 174698 592178 174934
rect 591942 139018 592178 139254
rect 591942 138698 592178 138934
rect 591942 103018 592178 103254
rect 591942 102698 592178 102934
rect 591942 67018 592178 67254
rect 591942 66698 592178 66934
rect 591942 31018 592178 31254
rect 591942 30698 592178 30934
rect 569786 -7022 570022 -6786
rect 569786 -7342 570022 -7106
rect 591942 -7022 592178 -6786
rect 591942 -7342 592178 -7106
<< metal5 >>
rect -8436 711300 -7836 711302
rect 29604 711300 30204 711302
rect 65604 711300 66204 711302
rect 101604 711300 102204 711302
rect 137604 711300 138204 711302
rect 173604 711300 174204 711302
rect 209604 711300 210204 711302
rect 245604 711300 246204 711302
rect 281604 711300 282204 711302
rect 317604 711300 318204 711302
rect 353604 711300 354204 711302
rect 389604 711300 390204 711302
rect 425604 711300 426204 711302
rect 461604 711300 462204 711302
rect 497604 711300 498204 711302
rect 533604 711300 534204 711302
rect 569604 711300 570204 711302
rect 591760 711300 592360 711302
rect -8436 711278 592360 711300
rect -8436 711042 -8254 711278
rect -8018 711042 29786 711278
rect 30022 711042 65786 711278
rect 66022 711042 101786 711278
rect 102022 711042 137786 711278
rect 138022 711042 173786 711278
rect 174022 711042 209786 711278
rect 210022 711042 245786 711278
rect 246022 711042 281786 711278
rect 282022 711042 317786 711278
rect 318022 711042 353786 711278
rect 354022 711042 389786 711278
rect 390022 711042 425786 711278
rect 426022 711042 461786 711278
rect 462022 711042 497786 711278
rect 498022 711042 533786 711278
rect 534022 711042 569786 711278
rect 570022 711042 591942 711278
rect 592178 711042 592360 711278
rect -8436 710958 592360 711042
rect -8436 710722 -8254 710958
rect -8018 710722 29786 710958
rect 30022 710722 65786 710958
rect 66022 710722 101786 710958
rect 102022 710722 137786 710958
rect 138022 710722 173786 710958
rect 174022 710722 209786 710958
rect 210022 710722 245786 710958
rect 246022 710722 281786 710958
rect 282022 710722 317786 710958
rect 318022 710722 353786 710958
rect 354022 710722 389786 710958
rect 390022 710722 425786 710958
rect 426022 710722 461786 710958
rect 462022 710722 497786 710958
rect 498022 710722 533786 710958
rect 534022 710722 569786 710958
rect 570022 710722 591942 710958
rect 592178 710722 592360 710958
rect -8436 710700 592360 710722
rect -8436 710698 -7836 710700
rect 29604 710698 30204 710700
rect 65604 710698 66204 710700
rect 101604 710698 102204 710700
rect 137604 710698 138204 710700
rect 173604 710698 174204 710700
rect 209604 710698 210204 710700
rect 245604 710698 246204 710700
rect 281604 710698 282204 710700
rect 317604 710698 318204 710700
rect 353604 710698 354204 710700
rect 389604 710698 390204 710700
rect 425604 710698 426204 710700
rect 461604 710698 462204 710700
rect 497604 710698 498204 710700
rect 533604 710698 534204 710700
rect 569604 710698 570204 710700
rect 591760 710698 592360 710700
rect -7516 710380 -6916 710382
rect 11604 710380 12204 710382
rect 47604 710380 48204 710382
rect 83604 710380 84204 710382
rect 119604 710380 120204 710382
rect 155604 710380 156204 710382
rect 191604 710380 192204 710382
rect 227604 710380 228204 710382
rect 263604 710380 264204 710382
rect 299604 710380 300204 710382
rect 335604 710380 336204 710382
rect 371604 710380 372204 710382
rect 407604 710380 408204 710382
rect 443604 710380 444204 710382
rect 479604 710380 480204 710382
rect 515604 710380 516204 710382
rect 551604 710380 552204 710382
rect 590840 710380 591440 710382
rect -7516 710358 591440 710380
rect -7516 710122 -7334 710358
rect -7098 710122 11786 710358
rect 12022 710122 47786 710358
rect 48022 710122 83786 710358
rect 84022 710122 119786 710358
rect 120022 710122 155786 710358
rect 156022 710122 191786 710358
rect 192022 710122 227786 710358
rect 228022 710122 263786 710358
rect 264022 710122 299786 710358
rect 300022 710122 335786 710358
rect 336022 710122 371786 710358
rect 372022 710122 407786 710358
rect 408022 710122 443786 710358
rect 444022 710122 479786 710358
rect 480022 710122 515786 710358
rect 516022 710122 551786 710358
rect 552022 710122 591022 710358
rect 591258 710122 591440 710358
rect -7516 710038 591440 710122
rect -7516 709802 -7334 710038
rect -7098 709802 11786 710038
rect 12022 709802 47786 710038
rect 48022 709802 83786 710038
rect 84022 709802 119786 710038
rect 120022 709802 155786 710038
rect 156022 709802 191786 710038
rect 192022 709802 227786 710038
rect 228022 709802 263786 710038
rect 264022 709802 299786 710038
rect 300022 709802 335786 710038
rect 336022 709802 371786 710038
rect 372022 709802 407786 710038
rect 408022 709802 443786 710038
rect 444022 709802 479786 710038
rect 480022 709802 515786 710038
rect 516022 709802 551786 710038
rect 552022 709802 591022 710038
rect 591258 709802 591440 710038
rect -7516 709780 591440 709802
rect -7516 709778 -6916 709780
rect 11604 709778 12204 709780
rect 47604 709778 48204 709780
rect 83604 709778 84204 709780
rect 119604 709778 120204 709780
rect 155604 709778 156204 709780
rect 191604 709778 192204 709780
rect 227604 709778 228204 709780
rect 263604 709778 264204 709780
rect 299604 709778 300204 709780
rect 335604 709778 336204 709780
rect 371604 709778 372204 709780
rect 407604 709778 408204 709780
rect 443604 709778 444204 709780
rect 479604 709778 480204 709780
rect 515604 709778 516204 709780
rect 551604 709778 552204 709780
rect 590840 709778 591440 709780
rect -6596 709460 -5996 709462
rect 26004 709460 26604 709462
rect 62004 709460 62604 709462
rect 98004 709460 98604 709462
rect 134004 709460 134604 709462
rect 170004 709460 170604 709462
rect 206004 709460 206604 709462
rect 242004 709460 242604 709462
rect 278004 709460 278604 709462
rect 314004 709460 314604 709462
rect 350004 709460 350604 709462
rect 386004 709460 386604 709462
rect 422004 709460 422604 709462
rect 458004 709460 458604 709462
rect 494004 709460 494604 709462
rect 530004 709460 530604 709462
rect 566004 709460 566604 709462
rect 589920 709460 590520 709462
rect -6596 709438 590520 709460
rect -6596 709202 -6414 709438
rect -6178 709202 26186 709438
rect 26422 709202 62186 709438
rect 62422 709202 98186 709438
rect 98422 709202 134186 709438
rect 134422 709202 170186 709438
rect 170422 709202 206186 709438
rect 206422 709202 242186 709438
rect 242422 709202 278186 709438
rect 278422 709202 314186 709438
rect 314422 709202 350186 709438
rect 350422 709202 386186 709438
rect 386422 709202 422186 709438
rect 422422 709202 458186 709438
rect 458422 709202 494186 709438
rect 494422 709202 530186 709438
rect 530422 709202 566186 709438
rect 566422 709202 590102 709438
rect 590338 709202 590520 709438
rect -6596 709118 590520 709202
rect -6596 708882 -6414 709118
rect -6178 708882 26186 709118
rect 26422 708882 62186 709118
rect 62422 708882 98186 709118
rect 98422 708882 134186 709118
rect 134422 708882 170186 709118
rect 170422 708882 206186 709118
rect 206422 708882 242186 709118
rect 242422 708882 278186 709118
rect 278422 708882 314186 709118
rect 314422 708882 350186 709118
rect 350422 708882 386186 709118
rect 386422 708882 422186 709118
rect 422422 708882 458186 709118
rect 458422 708882 494186 709118
rect 494422 708882 530186 709118
rect 530422 708882 566186 709118
rect 566422 708882 590102 709118
rect 590338 708882 590520 709118
rect -6596 708860 590520 708882
rect -6596 708858 -5996 708860
rect 26004 708858 26604 708860
rect 62004 708858 62604 708860
rect 98004 708858 98604 708860
rect 134004 708858 134604 708860
rect 170004 708858 170604 708860
rect 206004 708858 206604 708860
rect 242004 708858 242604 708860
rect 278004 708858 278604 708860
rect 314004 708858 314604 708860
rect 350004 708858 350604 708860
rect 386004 708858 386604 708860
rect 422004 708858 422604 708860
rect 458004 708858 458604 708860
rect 494004 708858 494604 708860
rect 530004 708858 530604 708860
rect 566004 708858 566604 708860
rect 589920 708858 590520 708860
rect -5676 708540 -5076 708542
rect 8004 708540 8604 708542
rect 44004 708540 44604 708542
rect 80004 708540 80604 708542
rect 116004 708540 116604 708542
rect 152004 708540 152604 708542
rect 188004 708540 188604 708542
rect 224004 708540 224604 708542
rect 260004 708540 260604 708542
rect 296004 708540 296604 708542
rect 332004 708540 332604 708542
rect 368004 708540 368604 708542
rect 404004 708540 404604 708542
rect 440004 708540 440604 708542
rect 476004 708540 476604 708542
rect 512004 708540 512604 708542
rect 548004 708540 548604 708542
rect 589000 708540 589600 708542
rect -5676 708518 589600 708540
rect -5676 708282 -5494 708518
rect -5258 708282 8186 708518
rect 8422 708282 44186 708518
rect 44422 708282 80186 708518
rect 80422 708282 116186 708518
rect 116422 708282 152186 708518
rect 152422 708282 188186 708518
rect 188422 708282 224186 708518
rect 224422 708282 260186 708518
rect 260422 708282 296186 708518
rect 296422 708282 332186 708518
rect 332422 708282 368186 708518
rect 368422 708282 404186 708518
rect 404422 708282 440186 708518
rect 440422 708282 476186 708518
rect 476422 708282 512186 708518
rect 512422 708282 548186 708518
rect 548422 708282 589182 708518
rect 589418 708282 589600 708518
rect -5676 708198 589600 708282
rect -5676 707962 -5494 708198
rect -5258 707962 8186 708198
rect 8422 707962 44186 708198
rect 44422 707962 80186 708198
rect 80422 707962 116186 708198
rect 116422 707962 152186 708198
rect 152422 707962 188186 708198
rect 188422 707962 224186 708198
rect 224422 707962 260186 708198
rect 260422 707962 296186 708198
rect 296422 707962 332186 708198
rect 332422 707962 368186 708198
rect 368422 707962 404186 708198
rect 404422 707962 440186 708198
rect 440422 707962 476186 708198
rect 476422 707962 512186 708198
rect 512422 707962 548186 708198
rect 548422 707962 589182 708198
rect 589418 707962 589600 708198
rect -5676 707940 589600 707962
rect -5676 707938 -5076 707940
rect 8004 707938 8604 707940
rect 44004 707938 44604 707940
rect 80004 707938 80604 707940
rect 116004 707938 116604 707940
rect 152004 707938 152604 707940
rect 188004 707938 188604 707940
rect 224004 707938 224604 707940
rect 260004 707938 260604 707940
rect 296004 707938 296604 707940
rect 332004 707938 332604 707940
rect 368004 707938 368604 707940
rect 404004 707938 404604 707940
rect 440004 707938 440604 707940
rect 476004 707938 476604 707940
rect 512004 707938 512604 707940
rect 548004 707938 548604 707940
rect 589000 707938 589600 707940
rect -4756 707620 -4156 707622
rect 22404 707620 23004 707622
rect 58404 707620 59004 707622
rect 94404 707620 95004 707622
rect 130404 707620 131004 707622
rect 166404 707620 167004 707622
rect 202404 707620 203004 707622
rect 238404 707620 239004 707622
rect 274404 707620 275004 707622
rect 310404 707620 311004 707622
rect 346404 707620 347004 707622
rect 382404 707620 383004 707622
rect 418404 707620 419004 707622
rect 454404 707620 455004 707622
rect 490404 707620 491004 707622
rect 526404 707620 527004 707622
rect 562404 707620 563004 707622
rect 588080 707620 588680 707622
rect -4756 707598 588680 707620
rect -4756 707362 -4574 707598
rect -4338 707362 22586 707598
rect 22822 707362 58586 707598
rect 58822 707362 94586 707598
rect 94822 707362 130586 707598
rect 130822 707362 166586 707598
rect 166822 707362 202586 707598
rect 202822 707362 238586 707598
rect 238822 707362 274586 707598
rect 274822 707362 310586 707598
rect 310822 707362 346586 707598
rect 346822 707362 382586 707598
rect 382822 707362 418586 707598
rect 418822 707362 454586 707598
rect 454822 707362 490586 707598
rect 490822 707362 526586 707598
rect 526822 707362 562586 707598
rect 562822 707362 588262 707598
rect 588498 707362 588680 707598
rect -4756 707278 588680 707362
rect -4756 707042 -4574 707278
rect -4338 707042 22586 707278
rect 22822 707042 58586 707278
rect 58822 707042 94586 707278
rect 94822 707042 130586 707278
rect 130822 707042 166586 707278
rect 166822 707042 202586 707278
rect 202822 707042 238586 707278
rect 238822 707042 274586 707278
rect 274822 707042 310586 707278
rect 310822 707042 346586 707278
rect 346822 707042 382586 707278
rect 382822 707042 418586 707278
rect 418822 707042 454586 707278
rect 454822 707042 490586 707278
rect 490822 707042 526586 707278
rect 526822 707042 562586 707278
rect 562822 707042 588262 707278
rect 588498 707042 588680 707278
rect -4756 707020 588680 707042
rect -4756 707018 -4156 707020
rect 22404 707018 23004 707020
rect 58404 707018 59004 707020
rect 94404 707018 95004 707020
rect 130404 707018 131004 707020
rect 166404 707018 167004 707020
rect 202404 707018 203004 707020
rect 238404 707018 239004 707020
rect 274404 707018 275004 707020
rect 310404 707018 311004 707020
rect 346404 707018 347004 707020
rect 382404 707018 383004 707020
rect 418404 707018 419004 707020
rect 454404 707018 455004 707020
rect 490404 707018 491004 707020
rect 526404 707018 527004 707020
rect 562404 707018 563004 707020
rect 588080 707018 588680 707020
rect -3836 706700 -3236 706702
rect 4404 706700 5004 706702
rect 40404 706700 41004 706702
rect 76404 706700 77004 706702
rect 112404 706700 113004 706702
rect 148404 706700 149004 706702
rect 184404 706700 185004 706702
rect 220404 706700 221004 706702
rect 256404 706700 257004 706702
rect 292404 706700 293004 706702
rect 328404 706700 329004 706702
rect 364404 706700 365004 706702
rect 400404 706700 401004 706702
rect 436404 706700 437004 706702
rect 472404 706700 473004 706702
rect 508404 706700 509004 706702
rect 544404 706700 545004 706702
rect 580404 706700 581004 706702
rect 587160 706700 587760 706702
rect -3836 706678 587760 706700
rect -3836 706442 -3654 706678
rect -3418 706442 4586 706678
rect 4822 706442 40586 706678
rect 40822 706442 76586 706678
rect 76822 706442 112586 706678
rect 112822 706442 148586 706678
rect 148822 706442 184586 706678
rect 184822 706442 220586 706678
rect 220822 706442 256586 706678
rect 256822 706442 292586 706678
rect 292822 706442 328586 706678
rect 328822 706442 364586 706678
rect 364822 706442 400586 706678
rect 400822 706442 436586 706678
rect 436822 706442 472586 706678
rect 472822 706442 508586 706678
rect 508822 706442 544586 706678
rect 544822 706442 580586 706678
rect 580822 706442 587342 706678
rect 587578 706442 587760 706678
rect -3836 706358 587760 706442
rect -3836 706122 -3654 706358
rect -3418 706122 4586 706358
rect 4822 706122 40586 706358
rect 40822 706122 76586 706358
rect 76822 706122 112586 706358
rect 112822 706122 148586 706358
rect 148822 706122 184586 706358
rect 184822 706122 220586 706358
rect 220822 706122 256586 706358
rect 256822 706122 292586 706358
rect 292822 706122 328586 706358
rect 328822 706122 364586 706358
rect 364822 706122 400586 706358
rect 400822 706122 436586 706358
rect 436822 706122 472586 706358
rect 472822 706122 508586 706358
rect 508822 706122 544586 706358
rect 544822 706122 580586 706358
rect 580822 706122 587342 706358
rect 587578 706122 587760 706358
rect -3836 706100 587760 706122
rect -3836 706098 -3236 706100
rect 4404 706098 5004 706100
rect 40404 706098 41004 706100
rect 76404 706098 77004 706100
rect 112404 706098 113004 706100
rect 148404 706098 149004 706100
rect 184404 706098 185004 706100
rect 220404 706098 221004 706100
rect 256404 706098 257004 706100
rect 292404 706098 293004 706100
rect 328404 706098 329004 706100
rect 364404 706098 365004 706100
rect 400404 706098 401004 706100
rect 436404 706098 437004 706100
rect 472404 706098 473004 706100
rect 508404 706098 509004 706100
rect 544404 706098 545004 706100
rect 580404 706098 581004 706100
rect 587160 706098 587760 706100
rect -2916 705780 -2316 705782
rect 18804 705780 19404 705782
rect 54804 705780 55404 705782
rect 90804 705780 91404 705782
rect 126804 705780 127404 705782
rect 162804 705780 163404 705782
rect 198804 705780 199404 705782
rect 234804 705780 235404 705782
rect 270804 705780 271404 705782
rect 306804 705780 307404 705782
rect 342804 705780 343404 705782
rect 378804 705780 379404 705782
rect 414804 705780 415404 705782
rect 450804 705780 451404 705782
rect 486804 705780 487404 705782
rect 522804 705780 523404 705782
rect 558804 705780 559404 705782
rect 586240 705780 586840 705782
rect -2916 705758 586840 705780
rect -2916 705522 -2734 705758
rect -2498 705522 18986 705758
rect 19222 705522 54986 705758
rect 55222 705522 90986 705758
rect 91222 705522 126986 705758
rect 127222 705522 162986 705758
rect 163222 705522 198986 705758
rect 199222 705522 234986 705758
rect 235222 705522 270986 705758
rect 271222 705522 306986 705758
rect 307222 705522 342986 705758
rect 343222 705522 378986 705758
rect 379222 705522 414986 705758
rect 415222 705522 450986 705758
rect 451222 705522 486986 705758
rect 487222 705522 522986 705758
rect 523222 705522 558986 705758
rect 559222 705522 586422 705758
rect 586658 705522 586840 705758
rect -2916 705438 586840 705522
rect -2916 705202 -2734 705438
rect -2498 705202 18986 705438
rect 19222 705202 54986 705438
rect 55222 705202 90986 705438
rect 91222 705202 126986 705438
rect 127222 705202 162986 705438
rect 163222 705202 198986 705438
rect 199222 705202 234986 705438
rect 235222 705202 270986 705438
rect 271222 705202 306986 705438
rect 307222 705202 342986 705438
rect 343222 705202 378986 705438
rect 379222 705202 414986 705438
rect 415222 705202 450986 705438
rect 451222 705202 486986 705438
rect 487222 705202 522986 705438
rect 523222 705202 558986 705438
rect 559222 705202 586422 705438
rect 586658 705202 586840 705438
rect -2916 705180 586840 705202
rect -2916 705178 -2316 705180
rect 18804 705178 19404 705180
rect 54804 705178 55404 705180
rect 90804 705178 91404 705180
rect 126804 705178 127404 705180
rect 162804 705178 163404 705180
rect 198804 705178 199404 705180
rect 234804 705178 235404 705180
rect 270804 705178 271404 705180
rect 306804 705178 307404 705180
rect 342804 705178 343404 705180
rect 378804 705178 379404 705180
rect 414804 705178 415404 705180
rect 450804 705178 451404 705180
rect 486804 705178 487404 705180
rect 522804 705178 523404 705180
rect 558804 705178 559404 705180
rect 586240 705178 586840 705180
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7516 697276 -6916 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590840 697276 591440 697278
rect -8436 697254 592360 697276
rect -8436 697018 -7334 697254
rect -7098 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591022 697254
rect 591258 697018 592360 697254
rect -8436 696934 592360 697018
rect -8436 696698 -7334 696934
rect -7098 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591022 696934
rect 591258 696698 592360 696934
rect -8436 696676 592360 696698
rect -7516 696674 -6916 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590840 696674 591440 696676
rect -5676 693676 -5076 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589000 693676 589600 693678
rect -6596 693654 590520 693676
rect -6596 693418 -5494 693654
rect -5258 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589182 693654
rect 589418 693418 590520 693654
rect -6596 693334 590520 693418
rect -6596 693098 -5494 693334
rect -5258 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589182 693334
rect 589418 693098 590520 693334
rect -6596 693076 590520 693098
rect -5676 693074 -5076 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589000 693074 589600 693076
rect -3836 690076 -3236 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587160 690076 587760 690078
rect -4756 690054 588680 690076
rect -4756 689818 -3654 690054
rect -3418 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587342 690054
rect 587578 689818 588680 690054
rect -4756 689734 588680 689818
rect -4756 689498 -3654 689734
rect -3418 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587342 689734
rect 587578 689498 588680 689734
rect -4756 689476 588680 689498
rect -3836 689474 -3236 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587160 689474 587760 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2916 686454 586840 686476
rect -2916 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586840 686454
rect -2916 686134 586840 686218
rect -2916 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586840 686134
rect -2916 685876 586840 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8436 679276 -7836 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591760 679276 592360 679278
rect -8436 679254 592360 679276
rect -8436 679018 -8254 679254
rect -8018 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 591942 679254
rect 592178 679018 592360 679254
rect -8436 678934 592360 679018
rect -8436 678698 -8254 678934
rect -8018 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 591942 678934
rect 592178 678698 592360 678934
rect -8436 678676 592360 678698
rect -8436 678674 -7836 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591760 678674 592360 678676
rect -6596 675676 -5996 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 589920 675676 590520 675678
rect -6596 675654 590520 675676
rect -6596 675418 -6414 675654
rect -6178 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590102 675654
rect 590338 675418 590520 675654
rect -6596 675334 590520 675418
rect -6596 675098 -6414 675334
rect -6178 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590102 675334
rect 590338 675098 590520 675334
rect -6596 675076 590520 675098
rect -6596 675074 -5996 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 589920 675074 590520 675076
rect -4756 672076 -4156 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588080 672076 588680 672078
rect -4756 672054 588680 672076
rect -4756 671818 -4574 672054
rect -4338 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588262 672054
rect 588498 671818 588680 672054
rect -4756 671734 588680 671818
rect -4756 671498 -4574 671734
rect -4338 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588262 671734
rect 588498 671498 588680 671734
rect -4756 671476 588680 671498
rect -4756 671474 -4156 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588080 671474 588680 671476
rect -2916 668476 -2316 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586240 668476 586840 668478
rect -2916 668454 586840 668476
rect -2916 668218 -2734 668454
rect -2498 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586422 668454
rect 586658 668218 586840 668454
rect -2916 668134 586840 668218
rect -2916 667898 -2734 668134
rect -2498 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586422 668134
rect 586658 667898 586840 668134
rect -2916 667876 586840 667898
rect -2916 667874 -2316 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586240 667874 586840 667876
rect -7516 661276 -6916 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590840 661276 591440 661278
rect -8436 661254 592360 661276
rect -8436 661018 -7334 661254
rect -7098 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591022 661254
rect 591258 661018 592360 661254
rect -8436 660934 592360 661018
rect -8436 660698 -7334 660934
rect -7098 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591022 660934
rect 591258 660698 592360 660934
rect -8436 660676 592360 660698
rect -7516 660674 -6916 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590840 660674 591440 660676
rect -5676 657676 -5076 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589000 657676 589600 657678
rect -6596 657654 590520 657676
rect -6596 657418 -5494 657654
rect -5258 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589182 657654
rect 589418 657418 590520 657654
rect -6596 657334 590520 657418
rect -6596 657098 -5494 657334
rect -5258 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589182 657334
rect 589418 657098 590520 657334
rect -6596 657076 590520 657098
rect -5676 657074 -5076 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589000 657074 589600 657076
rect -3836 654076 -3236 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587160 654076 587760 654078
rect -4756 654054 588680 654076
rect -4756 653818 -3654 654054
rect -3418 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587342 654054
rect 587578 653818 588680 654054
rect -4756 653734 588680 653818
rect -4756 653498 -3654 653734
rect -3418 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587342 653734
rect 587578 653498 588680 653734
rect -4756 653476 588680 653498
rect -3836 653474 -3236 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587160 653474 587760 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2916 650454 586840 650476
rect -2916 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586840 650454
rect -2916 650134 586840 650218
rect -2916 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586840 650134
rect -2916 649876 586840 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8436 643276 -7836 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 101604 643276 102204 643278
rect 137604 643276 138204 643278
rect 173604 643276 174204 643278
rect 209604 643276 210204 643278
rect 245604 643276 246204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591760 643276 592360 643278
rect -8436 643254 592360 643276
rect -8436 643018 -8254 643254
rect -8018 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 101786 643254
rect 102022 643018 137786 643254
rect 138022 643018 173786 643254
rect 174022 643018 209786 643254
rect 210022 643018 245786 643254
rect 246022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 591942 643254
rect 592178 643018 592360 643254
rect -8436 642934 592360 643018
rect -8436 642698 -8254 642934
rect -8018 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 101786 642934
rect 102022 642698 137786 642934
rect 138022 642698 173786 642934
rect 174022 642698 209786 642934
rect 210022 642698 245786 642934
rect 246022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 591942 642934
rect 592178 642698 592360 642934
rect -8436 642676 592360 642698
rect -8436 642674 -7836 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 101604 642674 102204 642676
rect 137604 642674 138204 642676
rect 173604 642674 174204 642676
rect 209604 642674 210204 642676
rect 245604 642674 246204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591760 642674 592360 642676
rect -6596 639676 -5996 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 98004 639676 98604 639678
rect 134004 639676 134604 639678
rect 170004 639676 170604 639678
rect 206004 639676 206604 639678
rect 242004 639676 242604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 589920 639676 590520 639678
rect -6596 639654 590520 639676
rect -6596 639418 -6414 639654
rect -6178 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 98186 639654
rect 98422 639418 134186 639654
rect 134422 639418 170186 639654
rect 170422 639418 206186 639654
rect 206422 639418 242186 639654
rect 242422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590102 639654
rect 590338 639418 590520 639654
rect -6596 639334 590520 639418
rect -6596 639098 -6414 639334
rect -6178 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 98186 639334
rect 98422 639098 134186 639334
rect 134422 639098 170186 639334
rect 170422 639098 206186 639334
rect 206422 639098 242186 639334
rect 242422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590102 639334
rect 590338 639098 590520 639334
rect -6596 639076 590520 639098
rect -6596 639074 -5996 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 98004 639074 98604 639076
rect 134004 639074 134604 639076
rect 170004 639074 170604 639076
rect 206004 639074 206604 639076
rect 242004 639074 242604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 589920 639074 590520 639076
rect -4756 636076 -4156 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588080 636076 588680 636078
rect -4756 636054 588680 636076
rect -4756 635818 -4574 636054
rect -4338 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588262 636054
rect 588498 635818 588680 636054
rect -4756 635734 588680 635818
rect -4756 635498 -4574 635734
rect -4338 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588262 635734
rect 588498 635498 588680 635734
rect -4756 635476 588680 635498
rect -4756 635474 -4156 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588080 635474 588680 635476
rect -2916 632476 -2316 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586240 632476 586840 632478
rect -2916 632454 586840 632476
rect -2916 632218 -2734 632454
rect -2498 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586422 632454
rect 586658 632218 586840 632454
rect -2916 632134 586840 632218
rect -2916 631898 -2734 632134
rect -2498 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586422 632134
rect 586658 631898 586840 632134
rect -2916 631876 586840 631898
rect -2916 631874 -2316 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586240 631874 586840 631876
rect -7516 625276 -6916 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 83604 625276 84204 625278
rect 119604 625276 120204 625278
rect 155604 625276 156204 625278
rect 191604 625276 192204 625278
rect 227604 625276 228204 625278
rect 263604 625276 264204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590840 625276 591440 625278
rect -8436 625254 592360 625276
rect -8436 625018 -7334 625254
rect -7098 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 83786 625254
rect 84022 625018 119786 625254
rect 120022 625018 155786 625254
rect 156022 625018 191786 625254
rect 192022 625018 227786 625254
rect 228022 625018 263786 625254
rect 264022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591022 625254
rect 591258 625018 592360 625254
rect -8436 624934 592360 625018
rect -8436 624698 -7334 624934
rect -7098 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 83786 624934
rect 84022 624698 119786 624934
rect 120022 624698 155786 624934
rect 156022 624698 191786 624934
rect 192022 624698 227786 624934
rect 228022 624698 263786 624934
rect 264022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591022 624934
rect 591258 624698 592360 624934
rect -8436 624676 592360 624698
rect -7516 624674 -6916 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 83604 624674 84204 624676
rect 119604 624674 120204 624676
rect 155604 624674 156204 624676
rect 191604 624674 192204 624676
rect 227604 624674 228204 624676
rect 263604 624674 264204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590840 624674 591440 624676
rect -5676 621676 -5076 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 80004 621676 80604 621678
rect 116004 621676 116604 621678
rect 152004 621676 152604 621678
rect 188004 621676 188604 621678
rect 224004 621676 224604 621678
rect 260004 621676 260604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589000 621676 589600 621678
rect -6596 621654 590520 621676
rect -6596 621418 -5494 621654
rect -5258 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 80186 621654
rect 80422 621418 116186 621654
rect 116422 621418 152186 621654
rect 152422 621418 188186 621654
rect 188422 621418 224186 621654
rect 224422 621418 260186 621654
rect 260422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589182 621654
rect 589418 621418 590520 621654
rect -6596 621334 590520 621418
rect -6596 621098 -5494 621334
rect -5258 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 80186 621334
rect 80422 621098 116186 621334
rect 116422 621098 152186 621334
rect 152422 621098 188186 621334
rect 188422 621098 224186 621334
rect 224422 621098 260186 621334
rect 260422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589182 621334
rect 589418 621098 590520 621334
rect -6596 621076 590520 621098
rect -5676 621074 -5076 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 80004 621074 80604 621076
rect 116004 621074 116604 621076
rect 152004 621074 152604 621076
rect 188004 621074 188604 621076
rect 224004 621074 224604 621076
rect 260004 621074 260604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589000 621074 589600 621076
rect -3836 618076 -3236 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587160 618076 587760 618078
rect -4756 618054 588680 618076
rect -4756 617818 -3654 618054
rect -3418 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587342 618054
rect 587578 617818 588680 618054
rect -4756 617734 588680 617818
rect -4756 617498 -3654 617734
rect -3418 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587342 617734
rect 587578 617498 588680 617734
rect -4756 617476 588680 617498
rect -3836 617474 -3236 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587160 617474 587760 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2916 614454 586840 614476
rect -2916 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586840 614454
rect -2916 614134 586840 614218
rect -2916 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586840 614134
rect -2916 613876 586840 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8436 607276 -7836 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 101604 607276 102204 607278
rect 137604 607276 138204 607278
rect 173604 607276 174204 607278
rect 209604 607276 210204 607278
rect 245604 607276 246204 607278
rect 281604 607276 282204 607278
rect 317604 607276 318204 607278
rect 353604 607276 354204 607278
rect 389604 607276 390204 607278
rect 425604 607276 426204 607278
rect 461604 607276 462204 607278
rect 497604 607276 498204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591760 607276 592360 607278
rect -8436 607254 592360 607276
rect -8436 607018 -8254 607254
rect -8018 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 101786 607254
rect 102022 607018 137786 607254
rect 138022 607018 173786 607254
rect 174022 607018 209786 607254
rect 210022 607018 245786 607254
rect 246022 607018 281786 607254
rect 282022 607018 317786 607254
rect 318022 607018 353786 607254
rect 354022 607018 389786 607254
rect 390022 607018 425786 607254
rect 426022 607018 461786 607254
rect 462022 607018 497786 607254
rect 498022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 591942 607254
rect 592178 607018 592360 607254
rect -8436 606934 592360 607018
rect -8436 606698 -8254 606934
rect -8018 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 101786 606934
rect 102022 606698 137786 606934
rect 138022 606698 173786 606934
rect 174022 606698 209786 606934
rect 210022 606698 245786 606934
rect 246022 606698 281786 606934
rect 282022 606698 317786 606934
rect 318022 606698 353786 606934
rect 354022 606698 389786 606934
rect 390022 606698 425786 606934
rect 426022 606698 461786 606934
rect 462022 606698 497786 606934
rect 498022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 591942 606934
rect 592178 606698 592360 606934
rect -8436 606676 592360 606698
rect -8436 606674 -7836 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 101604 606674 102204 606676
rect 137604 606674 138204 606676
rect 173604 606674 174204 606676
rect 209604 606674 210204 606676
rect 245604 606674 246204 606676
rect 281604 606674 282204 606676
rect 317604 606674 318204 606676
rect 353604 606674 354204 606676
rect 389604 606674 390204 606676
rect 425604 606674 426204 606676
rect 461604 606674 462204 606676
rect 497604 606674 498204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591760 606674 592360 606676
rect -6596 603676 -5996 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 98004 603676 98604 603678
rect 134004 603676 134604 603678
rect 170004 603676 170604 603678
rect 206004 603676 206604 603678
rect 242004 603676 242604 603678
rect 278004 603676 278604 603678
rect 314004 603676 314604 603678
rect 350004 603676 350604 603678
rect 386004 603676 386604 603678
rect 422004 603676 422604 603678
rect 458004 603676 458604 603678
rect 494004 603676 494604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 589920 603676 590520 603678
rect -6596 603654 590520 603676
rect -6596 603418 -6414 603654
rect -6178 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 98186 603654
rect 98422 603418 134186 603654
rect 134422 603418 170186 603654
rect 170422 603418 206186 603654
rect 206422 603418 242186 603654
rect 242422 603418 278186 603654
rect 278422 603418 314186 603654
rect 314422 603418 350186 603654
rect 350422 603418 386186 603654
rect 386422 603418 422186 603654
rect 422422 603418 458186 603654
rect 458422 603418 494186 603654
rect 494422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590102 603654
rect 590338 603418 590520 603654
rect -6596 603334 590520 603418
rect -6596 603098 -6414 603334
rect -6178 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 98186 603334
rect 98422 603098 134186 603334
rect 134422 603098 170186 603334
rect 170422 603098 206186 603334
rect 206422 603098 242186 603334
rect 242422 603098 278186 603334
rect 278422 603098 314186 603334
rect 314422 603098 350186 603334
rect 350422 603098 386186 603334
rect 386422 603098 422186 603334
rect 422422 603098 458186 603334
rect 458422 603098 494186 603334
rect 494422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590102 603334
rect 590338 603098 590520 603334
rect -6596 603076 590520 603098
rect -6596 603074 -5996 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 98004 603074 98604 603076
rect 134004 603074 134604 603076
rect 170004 603074 170604 603076
rect 206004 603074 206604 603076
rect 242004 603074 242604 603076
rect 278004 603074 278604 603076
rect 314004 603074 314604 603076
rect 350004 603074 350604 603076
rect 386004 603074 386604 603076
rect 422004 603074 422604 603076
rect 458004 603074 458604 603076
rect 494004 603074 494604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 589920 603074 590520 603076
rect -4756 600076 -4156 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 94404 600076 95004 600078
rect 130404 600076 131004 600078
rect 166404 600076 167004 600078
rect 202404 600076 203004 600078
rect 238404 600076 239004 600078
rect 274404 600076 275004 600078
rect 310404 600076 311004 600078
rect 346404 600076 347004 600078
rect 382404 600076 383004 600078
rect 418404 600076 419004 600078
rect 454404 600076 455004 600078
rect 490404 600076 491004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588080 600076 588680 600078
rect -4756 600054 588680 600076
rect -4756 599818 -4574 600054
rect -4338 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 94586 600054
rect 94822 599818 130586 600054
rect 130822 599818 166586 600054
rect 166822 599818 202586 600054
rect 202822 599818 238586 600054
rect 238822 599818 274586 600054
rect 274822 599818 310586 600054
rect 310822 599818 346586 600054
rect 346822 599818 382586 600054
rect 382822 599818 418586 600054
rect 418822 599818 454586 600054
rect 454822 599818 490586 600054
rect 490822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588262 600054
rect 588498 599818 588680 600054
rect -4756 599734 588680 599818
rect -4756 599498 -4574 599734
rect -4338 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 94586 599734
rect 94822 599498 130586 599734
rect 130822 599498 166586 599734
rect 166822 599498 202586 599734
rect 202822 599498 238586 599734
rect 238822 599498 274586 599734
rect 274822 599498 310586 599734
rect 310822 599498 346586 599734
rect 346822 599498 382586 599734
rect 382822 599498 418586 599734
rect 418822 599498 454586 599734
rect 454822 599498 490586 599734
rect 490822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588262 599734
rect 588498 599498 588680 599734
rect -4756 599476 588680 599498
rect -4756 599474 -4156 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 94404 599474 95004 599476
rect 130404 599474 131004 599476
rect 166404 599474 167004 599476
rect 202404 599474 203004 599476
rect 238404 599474 239004 599476
rect 274404 599474 275004 599476
rect 310404 599474 311004 599476
rect 346404 599474 347004 599476
rect 382404 599474 383004 599476
rect 418404 599474 419004 599476
rect 454404 599474 455004 599476
rect 490404 599474 491004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588080 599474 588680 599476
rect -2916 596476 -2316 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586240 596476 586840 596478
rect -2916 596454 586840 596476
rect -2916 596218 -2734 596454
rect -2498 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586422 596454
rect 586658 596218 586840 596454
rect -2916 596134 586840 596218
rect -2916 595898 -2734 596134
rect -2498 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586422 596134
rect 586658 595898 586840 596134
rect -2916 595876 586840 595898
rect -2916 595874 -2316 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586240 595874 586840 595876
rect -7516 589276 -6916 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 83604 589276 84204 589278
rect 119604 589276 120204 589278
rect 155604 589276 156204 589278
rect 191604 589276 192204 589278
rect 227604 589276 228204 589278
rect 263604 589276 264204 589278
rect 299604 589276 300204 589278
rect 335604 589276 336204 589278
rect 371604 589276 372204 589278
rect 407604 589276 408204 589278
rect 443604 589276 444204 589278
rect 479604 589276 480204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590840 589276 591440 589278
rect -8436 589254 592360 589276
rect -8436 589018 -7334 589254
rect -7098 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 83786 589254
rect 84022 589018 119786 589254
rect 120022 589018 155786 589254
rect 156022 589018 191786 589254
rect 192022 589018 227786 589254
rect 228022 589018 263786 589254
rect 264022 589018 299786 589254
rect 300022 589018 335786 589254
rect 336022 589018 371786 589254
rect 372022 589018 407786 589254
rect 408022 589018 443786 589254
rect 444022 589018 479786 589254
rect 480022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591022 589254
rect 591258 589018 592360 589254
rect -8436 588934 592360 589018
rect -8436 588698 -7334 588934
rect -7098 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 83786 588934
rect 84022 588698 119786 588934
rect 120022 588698 155786 588934
rect 156022 588698 191786 588934
rect 192022 588698 227786 588934
rect 228022 588698 263786 588934
rect 264022 588698 299786 588934
rect 300022 588698 335786 588934
rect 336022 588698 371786 588934
rect 372022 588698 407786 588934
rect 408022 588698 443786 588934
rect 444022 588698 479786 588934
rect 480022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591022 588934
rect 591258 588698 592360 588934
rect -8436 588676 592360 588698
rect -7516 588674 -6916 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 83604 588674 84204 588676
rect 119604 588674 120204 588676
rect 155604 588674 156204 588676
rect 191604 588674 192204 588676
rect 227604 588674 228204 588676
rect 263604 588674 264204 588676
rect 299604 588674 300204 588676
rect 335604 588674 336204 588676
rect 371604 588674 372204 588676
rect 407604 588674 408204 588676
rect 443604 588674 444204 588676
rect 479604 588674 480204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590840 588674 591440 588676
rect -5676 585676 -5076 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 80004 585676 80604 585678
rect 116004 585676 116604 585678
rect 152004 585676 152604 585678
rect 188004 585676 188604 585678
rect 224004 585676 224604 585678
rect 260004 585676 260604 585678
rect 296004 585676 296604 585678
rect 332004 585676 332604 585678
rect 368004 585676 368604 585678
rect 404004 585676 404604 585678
rect 440004 585676 440604 585678
rect 476004 585676 476604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589000 585676 589600 585678
rect -6596 585654 590520 585676
rect -6596 585418 -5494 585654
rect -5258 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 80186 585654
rect 80422 585418 116186 585654
rect 116422 585418 152186 585654
rect 152422 585418 188186 585654
rect 188422 585418 224186 585654
rect 224422 585418 260186 585654
rect 260422 585418 296186 585654
rect 296422 585418 332186 585654
rect 332422 585418 368186 585654
rect 368422 585418 404186 585654
rect 404422 585418 440186 585654
rect 440422 585418 476186 585654
rect 476422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589182 585654
rect 589418 585418 590520 585654
rect -6596 585334 590520 585418
rect -6596 585098 -5494 585334
rect -5258 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 80186 585334
rect 80422 585098 116186 585334
rect 116422 585098 152186 585334
rect 152422 585098 188186 585334
rect 188422 585098 224186 585334
rect 224422 585098 260186 585334
rect 260422 585098 296186 585334
rect 296422 585098 332186 585334
rect 332422 585098 368186 585334
rect 368422 585098 404186 585334
rect 404422 585098 440186 585334
rect 440422 585098 476186 585334
rect 476422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589182 585334
rect 589418 585098 590520 585334
rect -6596 585076 590520 585098
rect -5676 585074 -5076 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 80004 585074 80604 585076
rect 116004 585074 116604 585076
rect 152004 585074 152604 585076
rect 188004 585074 188604 585076
rect 224004 585074 224604 585076
rect 260004 585074 260604 585076
rect 296004 585074 296604 585076
rect 332004 585074 332604 585076
rect 368004 585074 368604 585076
rect 404004 585074 404604 585076
rect 440004 585074 440604 585076
rect 476004 585074 476604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589000 585074 589600 585076
rect -3836 582076 -3236 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 112404 582076 113004 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 220404 582076 221004 582078
rect 256404 582076 257004 582078
rect 292404 582076 293004 582078
rect 328404 582076 329004 582078
rect 364404 582076 365004 582078
rect 400404 582076 401004 582078
rect 436404 582076 437004 582078
rect 472404 582076 473004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587160 582076 587760 582078
rect -4756 582054 588680 582076
rect -4756 581818 -3654 582054
rect -3418 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 112586 582054
rect 112822 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 220586 582054
rect 220822 581818 256586 582054
rect 256822 581818 292586 582054
rect 292822 581818 328586 582054
rect 328822 581818 364586 582054
rect 364822 581818 400586 582054
rect 400822 581818 436586 582054
rect 436822 581818 472586 582054
rect 472822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587342 582054
rect 587578 581818 588680 582054
rect -4756 581734 588680 581818
rect -4756 581498 -3654 581734
rect -3418 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 112586 581734
rect 112822 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 220586 581734
rect 220822 581498 256586 581734
rect 256822 581498 292586 581734
rect 292822 581498 328586 581734
rect 328822 581498 364586 581734
rect 364822 581498 400586 581734
rect 400822 581498 436586 581734
rect 436822 581498 472586 581734
rect 472822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587342 581734
rect 587578 581498 588680 581734
rect -4756 581476 588680 581498
rect -3836 581474 -3236 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 112404 581474 113004 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 220404 581474 221004 581476
rect 256404 581474 257004 581476
rect 292404 581474 293004 581476
rect 328404 581474 329004 581476
rect 364404 581474 365004 581476
rect 400404 581474 401004 581476
rect 436404 581474 437004 581476
rect 472404 581474 473004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587160 581474 587760 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 108804 578476 109404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 216804 578476 217404 578478
rect 252804 578476 253404 578478
rect 288804 578476 289404 578478
rect 324804 578476 325404 578478
rect 360804 578476 361404 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 468804 578476 469404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2916 578454 586840 578476
rect -2916 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 324986 578454
rect 325222 578218 360986 578454
rect 361222 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586840 578454
rect -2916 578134 586840 578218
rect -2916 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 324986 578134
rect 325222 577898 360986 578134
rect 361222 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586840 578134
rect -2916 577876 586840 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 108804 577874 109404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 216804 577874 217404 577876
rect 252804 577874 253404 577876
rect 288804 577874 289404 577876
rect 324804 577874 325404 577876
rect 360804 577874 361404 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 468804 577874 469404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8436 571276 -7836 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 101604 571276 102204 571278
rect 137604 571276 138204 571278
rect 173604 571276 174204 571278
rect 209604 571276 210204 571278
rect 245604 571276 246204 571278
rect 281604 571276 282204 571278
rect 317604 571276 318204 571278
rect 353604 571276 354204 571278
rect 389604 571276 390204 571278
rect 425604 571276 426204 571278
rect 461604 571276 462204 571278
rect 497604 571276 498204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591760 571276 592360 571278
rect -8436 571254 592360 571276
rect -8436 571018 -8254 571254
rect -8018 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 101786 571254
rect 102022 571018 137786 571254
rect 138022 571018 173786 571254
rect 174022 571018 209786 571254
rect 210022 571018 245786 571254
rect 246022 571018 281786 571254
rect 282022 571018 317786 571254
rect 318022 571018 353786 571254
rect 354022 571018 389786 571254
rect 390022 571018 425786 571254
rect 426022 571018 461786 571254
rect 462022 571018 497786 571254
rect 498022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 591942 571254
rect 592178 571018 592360 571254
rect -8436 570934 592360 571018
rect -8436 570698 -8254 570934
rect -8018 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 101786 570934
rect 102022 570698 137786 570934
rect 138022 570698 173786 570934
rect 174022 570698 209786 570934
rect 210022 570698 245786 570934
rect 246022 570698 281786 570934
rect 282022 570698 317786 570934
rect 318022 570698 353786 570934
rect 354022 570698 389786 570934
rect 390022 570698 425786 570934
rect 426022 570698 461786 570934
rect 462022 570698 497786 570934
rect 498022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 591942 570934
rect 592178 570698 592360 570934
rect -8436 570676 592360 570698
rect -8436 570674 -7836 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 101604 570674 102204 570676
rect 137604 570674 138204 570676
rect 173604 570674 174204 570676
rect 209604 570674 210204 570676
rect 245604 570674 246204 570676
rect 281604 570674 282204 570676
rect 317604 570674 318204 570676
rect 353604 570674 354204 570676
rect 389604 570674 390204 570676
rect 425604 570674 426204 570676
rect 461604 570674 462204 570676
rect 497604 570674 498204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591760 570674 592360 570676
rect -6596 567676 -5996 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 98004 567676 98604 567678
rect 134004 567676 134604 567678
rect 170004 567676 170604 567678
rect 206004 567676 206604 567678
rect 242004 567676 242604 567678
rect 278004 567676 278604 567678
rect 314004 567676 314604 567678
rect 350004 567676 350604 567678
rect 386004 567676 386604 567678
rect 422004 567676 422604 567678
rect 458004 567676 458604 567678
rect 494004 567676 494604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 589920 567676 590520 567678
rect -6596 567654 590520 567676
rect -6596 567418 -6414 567654
rect -6178 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 98186 567654
rect 98422 567418 134186 567654
rect 134422 567418 170186 567654
rect 170422 567418 206186 567654
rect 206422 567418 242186 567654
rect 242422 567418 278186 567654
rect 278422 567418 314186 567654
rect 314422 567418 350186 567654
rect 350422 567418 386186 567654
rect 386422 567418 422186 567654
rect 422422 567418 458186 567654
rect 458422 567418 494186 567654
rect 494422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590102 567654
rect 590338 567418 590520 567654
rect -6596 567334 590520 567418
rect -6596 567098 -6414 567334
rect -6178 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 98186 567334
rect 98422 567098 134186 567334
rect 134422 567098 170186 567334
rect 170422 567098 206186 567334
rect 206422 567098 242186 567334
rect 242422 567098 278186 567334
rect 278422 567098 314186 567334
rect 314422 567098 350186 567334
rect 350422 567098 386186 567334
rect 386422 567098 422186 567334
rect 422422 567098 458186 567334
rect 458422 567098 494186 567334
rect 494422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590102 567334
rect 590338 567098 590520 567334
rect -6596 567076 590520 567098
rect -6596 567074 -5996 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 98004 567074 98604 567076
rect 134004 567074 134604 567076
rect 170004 567074 170604 567076
rect 206004 567074 206604 567076
rect 242004 567074 242604 567076
rect 278004 567074 278604 567076
rect 314004 567074 314604 567076
rect 350004 567074 350604 567076
rect 386004 567074 386604 567076
rect 422004 567074 422604 567076
rect 458004 567074 458604 567076
rect 494004 567074 494604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 589920 567074 590520 567076
rect -4756 564076 -4156 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 94404 564076 95004 564078
rect 130404 564076 131004 564078
rect 166404 564076 167004 564078
rect 202404 564076 203004 564078
rect 238404 564076 239004 564078
rect 274404 564076 275004 564078
rect 310404 564076 311004 564078
rect 346404 564076 347004 564078
rect 382404 564076 383004 564078
rect 418404 564076 419004 564078
rect 454404 564076 455004 564078
rect 490404 564076 491004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588080 564076 588680 564078
rect -4756 564054 588680 564076
rect -4756 563818 -4574 564054
rect -4338 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 94586 564054
rect 94822 563818 130586 564054
rect 130822 563818 166586 564054
rect 166822 563818 202586 564054
rect 202822 563818 238586 564054
rect 238822 563818 274586 564054
rect 274822 563818 310586 564054
rect 310822 563818 346586 564054
rect 346822 563818 382586 564054
rect 382822 563818 418586 564054
rect 418822 563818 454586 564054
rect 454822 563818 490586 564054
rect 490822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588262 564054
rect 588498 563818 588680 564054
rect -4756 563734 588680 563818
rect -4756 563498 -4574 563734
rect -4338 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 94586 563734
rect 94822 563498 130586 563734
rect 130822 563498 166586 563734
rect 166822 563498 202586 563734
rect 202822 563498 238586 563734
rect 238822 563498 274586 563734
rect 274822 563498 310586 563734
rect 310822 563498 346586 563734
rect 346822 563498 382586 563734
rect 382822 563498 418586 563734
rect 418822 563498 454586 563734
rect 454822 563498 490586 563734
rect 490822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588262 563734
rect 588498 563498 588680 563734
rect -4756 563476 588680 563498
rect -4756 563474 -4156 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 94404 563474 95004 563476
rect 130404 563474 131004 563476
rect 166404 563474 167004 563476
rect 202404 563474 203004 563476
rect 238404 563474 239004 563476
rect 274404 563474 275004 563476
rect 310404 563474 311004 563476
rect 346404 563474 347004 563476
rect 382404 563474 383004 563476
rect 418404 563474 419004 563476
rect 454404 563474 455004 563476
rect 490404 563474 491004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588080 563474 588680 563476
rect -2916 560476 -2316 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 342804 560476 343404 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586240 560476 586840 560478
rect -2916 560454 586840 560476
rect -2916 560218 -2734 560454
rect -2498 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 342986 560454
rect 343222 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586422 560454
rect 586658 560218 586840 560454
rect -2916 560134 586840 560218
rect -2916 559898 -2734 560134
rect -2498 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 342986 560134
rect 343222 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586422 560134
rect 586658 559898 586840 560134
rect -2916 559876 586840 559898
rect -2916 559874 -2316 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 342804 559874 343404 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586240 559874 586840 559876
rect -7516 553276 -6916 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 83604 553276 84204 553278
rect 119604 553276 120204 553278
rect 155604 553276 156204 553278
rect 191604 553276 192204 553278
rect 227604 553276 228204 553278
rect 263604 553276 264204 553278
rect 299604 553276 300204 553278
rect 335604 553276 336204 553278
rect 371604 553276 372204 553278
rect 407604 553276 408204 553278
rect 443604 553276 444204 553278
rect 479604 553276 480204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590840 553276 591440 553278
rect -8436 553254 592360 553276
rect -8436 553018 -7334 553254
rect -7098 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 83786 553254
rect 84022 553018 119786 553254
rect 120022 553018 155786 553254
rect 156022 553018 191786 553254
rect 192022 553018 227786 553254
rect 228022 553018 263786 553254
rect 264022 553018 299786 553254
rect 300022 553018 335786 553254
rect 336022 553018 371786 553254
rect 372022 553018 407786 553254
rect 408022 553018 443786 553254
rect 444022 553018 479786 553254
rect 480022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591022 553254
rect 591258 553018 592360 553254
rect -8436 552934 592360 553018
rect -8436 552698 -7334 552934
rect -7098 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 83786 552934
rect 84022 552698 119786 552934
rect 120022 552698 155786 552934
rect 156022 552698 191786 552934
rect 192022 552698 227786 552934
rect 228022 552698 263786 552934
rect 264022 552698 299786 552934
rect 300022 552698 335786 552934
rect 336022 552698 371786 552934
rect 372022 552698 407786 552934
rect 408022 552698 443786 552934
rect 444022 552698 479786 552934
rect 480022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591022 552934
rect 591258 552698 592360 552934
rect -8436 552676 592360 552698
rect -7516 552674 -6916 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 83604 552674 84204 552676
rect 119604 552674 120204 552676
rect 155604 552674 156204 552676
rect 191604 552674 192204 552676
rect 227604 552674 228204 552676
rect 263604 552674 264204 552676
rect 299604 552674 300204 552676
rect 335604 552674 336204 552676
rect 371604 552674 372204 552676
rect 407604 552674 408204 552676
rect 443604 552674 444204 552676
rect 479604 552674 480204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590840 552674 591440 552676
rect -5676 549676 -5076 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 116004 549676 116604 549678
rect 152004 549676 152604 549678
rect 188004 549676 188604 549678
rect 224004 549676 224604 549678
rect 260004 549676 260604 549678
rect 296004 549676 296604 549678
rect 332004 549676 332604 549678
rect 368004 549676 368604 549678
rect 404004 549676 404604 549678
rect 440004 549676 440604 549678
rect 476004 549676 476604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589000 549676 589600 549678
rect -6596 549654 590520 549676
rect -6596 549418 -5494 549654
rect -5258 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 116186 549654
rect 116422 549418 152186 549654
rect 152422 549418 188186 549654
rect 188422 549418 224186 549654
rect 224422 549418 260186 549654
rect 260422 549418 296186 549654
rect 296422 549418 332186 549654
rect 332422 549418 368186 549654
rect 368422 549418 404186 549654
rect 404422 549418 440186 549654
rect 440422 549418 476186 549654
rect 476422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589182 549654
rect 589418 549418 590520 549654
rect -6596 549334 590520 549418
rect -6596 549098 -5494 549334
rect -5258 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 116186 549334
rect 116422 549098 152186 549334
rect 152422 549098 188186 549334
rect 188422 549098 224186 549334
rect 224422 549098 260186 549334
rect 260422 549098 296186 549334
rect 296422 549098 332186 549334
rect 332422 549098 368186 549334
rect 368422 549098 404186 549334
rect 404422 549098 440186 549334
rect 440422 549098 476186 549334
rect 476422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589182 549334
rect 589418 549098 590520 549334
rect -6596 549076 590520 549098
rect -5676 549074 -5076 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 116004 549074 116604 549076
rect 152004 549074 152604 549076
rect 188004 549074 188604 549076
rect 224004 549074 224604 549076
rect 260004 549074 260604 549076
rect 296004 549074 296604 549076
rect 332004 549074 332604 549076
rect 368004 549074 368604 549076
rect 404004 549074 404604 549076
rect 440004 549074 440604 549076
rect 476004 549074 476604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589000 549074 589600 549076
rect -3836 546076 -3236 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 112404 546076 113004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 328404 546076 329004 546078
rect 364404 546076 365004 546078
rect 400404 546076 401004 546078
rect 436404 546076 437004 546078
rect 472404 546076 473004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587160 546076 587760 546078
rect -4756 546054 588680 546076
rect -4756 545818 -3654 546054
rect -3418 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 112586 546054
rect 112822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 328586 546054
rect 328822 545818 364586 546054
rect 364822 545818 400586 546054
rect 400822 545818 436586 546054
rect 436822 545818 472586 546054
rect 472822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587342 546054
rect 587578 545818 588680 546054
rect -4756 545734 588680 545818
rect -4756 545498 -3654 545734
rect -3418 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 112586 545734
rect 112822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 328586 545734
rect 328822 545498 364586 545734
rect 364822 545498 400586 545734
rect 400822 545498 436586 545734
rect 436822 545498 472586 545734
rect 472822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587342 545734
rect 587578 545498 588680 545734
rect -4756 545476 588680 545498
rect -3836 545474 -3236 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 112404 545474 113004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 328404 545474 329004 545476
rect 364404 545474 365004 545476
rect 400404 545474 401004 545476
rect 436404 545474 437004 545476
rect 472404 545474 473004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587160 545474 587760 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 108804 542476 109404 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 216804 542476 217404 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2916 542454 586840 542476
rect -2916 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 216986 542454
rect 217222 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586840 542454
rect -2916 542134 586840 542218
rect -2916 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 216986 542134
rect 217222 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586840 542134
rect -2916 541876 586840 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 108804 541874 109404 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 216804 541874 217404 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8436 535276 -7836 535278
rect 29604 535276 30204 535278
rect 65604 535276 66204 535278
rect 101604 535276 102204 535278
rect 137604 535276 138204 535278
rect 173604 535276 174204 535278
rect 209604 535276 210204 535278
rect 245604 535276 246204 535278
rect 281604 535276 282204 535278
rect 317604 535276 318204 535278
rect 353604 535276 354204 535278
rect 389604 535276 390204 535278
rect 425604 535276 426204 535278
rect 461604 535276 462204 535278
rect 497604 535276 498204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591760 535276 592360 535278
rect -8436 535254 592360 535276
rect -8436 535018 -8254 535254
rect -8018 535018 29786 535254
rect 30022 535018 65786 535254
rect 66022 535018 101786 535254
rect 102022 535018 137786 535254
rect 138022 535018 173786 535254
rect 174022 535018 209786 535254
rect 210022 535018 245786 535254
rect 246022 535018 281786 535254
rect 282022 535018 317786 535254
rect 318022 535018 353786 535254
rect 354022 535018 389786 535254
rect 390022 535018 425786 535254
rect 426022 535018 461786 535254
rect 462022 535018 497786 535254
rect 498022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 591942 535254
rect 592178 535018 592360 535254
rect -8436 534934 592360 535018
rect -8436 534698 -8254 534934
rect -8018 534698 29786 534934
rect 30022 534698 65786 534934
rect 66022 534698 101786 534934
rect 102022 534698 137786 534934
rect 138022 534698 173786 534934
rect 174022 534698 209786 534934
rect 210022 534698 245786 534934
rect 246022 534698 281786 534934
rect 282022 534698 317786 534934
rect 318022 534698 353786 534934
rect 354022 534698 389786 534934
rect 390022 534698 425786 534934
rect 426022 534698 461786 534934
rect 462022 534698 497786 534934
rect 498022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 591942 534934
rect 592178 534698 592360 534934
rect -8436 534676 592360 534698
rect -8436 534674 -7836 534676
rect 29604 534674 30204 534676
rect 65604 534674 66204 534676
rect 101604 534674 102204 534676
rect 137604 534674 138204 534676
rect 173604 534674 174204 534676
rect 209604 534674 210204 534676
rect 245604 534674 246204 534676
rect 281604 534674 282204 534676
rect 317604 534674 318204 534676
rect 353604 534674 354204 534676
rect 389604 534674 390204 534676
rect 425604 534674 426204 534676
rect 461604 534674 462204 534676
rect 497604 534674 498204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591760 534674 592360 534676
rect -6596 531676 -5996 531678
rect 26004 531676 26604 531678
rect 62004 531676 62604 531678
rect 98004 531676 98604 531678
rect 134004 531676 134604 531678
rect 170004 531676 170604 531678
rect 206004 531676 206604 531678
rect 242004 531676 242604 531678
rect 278004 531676 278604 531678
rect 314004 531676 314604 531678
rect 350004 531676 350604 531678
rect 386004 531676 386604 531678
rect 422004 531676 422604 531678
rect 458004 531676 458604 531678
rect 494004 531676 494604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 589920 531676 590520 531678
rect -6596 531654 590520 531676
rect -6596 531418 -6414 531654
rect -6178 531418 26186 531654
rect 26422 531418 62186 531654
rect 62422 531418 98186 531654
rect 98422 531418 134186 531654
rect 134422 531418 170186 531654
rect 170422 531418 206186 531654
rect 206422 531418 242186 531654
rect 242422 531418 278186 531654
rect 278422 531418 314186 531654
rect 314422 531418 350186 531654
rect 350422 531418 386186 531654
rect 386422 531418 422186 531654
rect 422422 531418 458186 531654
rect 458422 531418 494186 531654
rect 494422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590102 531654
rect 590338 531418 590520 531654
rect -6596 531334 590520 531418
rect -6596 531098 -6414 531334
rect -6178 531098 26186 531334
rect 26422 531098 62186 531334
rect 62422 531098 98186 531334
rect 98422 531098 134186 531334
rect 134422 531098 170186 531334
rect 170422 531098 206186 531334
rect 206422 531098 242186 531334
rect 242422 531098 278186 531334
rect 278422 531098 314186 531334
rect 314422 531098 350186 531334
rect 350422 531098 386186 531334
rect 386422 531098 422186 531334
rect 422422 531098 458186 531334
rect 458422 531098 494186 531334
rect 494422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590102 531334
rect 590338 531098 590520 531334
rect -6596 531076 590520 531098
rect -6596 531074 -5996 531076
rect 26004 531074 26604 531076
rect 62004 531074 62604 531076
rect 98004 531074 98604 531076
rect 134004 531074 134604 531076
rect 170004 531074 170604 531076
rect 206004 531074 206604 531076
rect 242004 531074 242604 531076
rect 278004 531074 278604 531076
rect 314004 531074 314604 531076
rect 350004 531074 350604 531076
rect 386004 531074 386604 531076
rect 422004 531074 422604 531076
rect 458004 531074 458604 531076
rect 494004 531074 494604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 589920 531074 590520 531076
rect -4756 528076 -4156 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 94404 528076 95004 528078
rect 130404 528076 131004 528078
rect 166404 528076 167004 528078
rect 202404 528076 203004 528078
rect 238404 528076 239004 528078
rect 274404 528076 275004 528078
rect 310404 528076 311004 528078
rect 346404 528076 347004 528078
rect 382404 528076 383004 528078
rect 418404 528076 419004 528078
rect 454404 528076 455004 528078
rect 490404 528076 491004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588080 528076 588680 528078
rect -4756 528054 588680 528076
rect -4756 527818 -4574 528054
rect -4338 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 94586 528054
rect 94822 527818 130586 528054
rect 130822 527818 166586 528054
rect 166822 527818 202586 528054
rect 202822 527818 238586 528054
rect 238822 527818 274586 528054
rect 274822 527818 310586 528054
rect 310822 527818 346586 528054
rect 346822 527818 382586 528054
rect 382822 527818 418586 528054
rect 418822 527818 454586 528054
rect 454822 527818 490586 528054
rect 490822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588262 528054
rect 588498 527818 588680 528054
rect -4756 527734 588680 527818
rect -4756 527498 -4574 527734
rect -4338 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 94586 527734
rect 94822 527498 130586 527734
rect 130822 527498 166586 527734
rect 166822 527498 202586 527734
rect 202822 527498 238586 527734
rect 238822 527498 274586 527734
rect 274822 527498 310586 527734
rect 310822 527498 346586 527734
rect 346822 527498 382586 527734
rect 382822 527498 418586 527734
rect 418822 527498 454586 527734
rect 454822 527498 490586 527734
rect 490822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588262 527734
rect 588498 527498 588680 527734
rect -4756 527476 588680 527498
rect -4756 527474 -4156 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 94404 527474 95004 527476
rect 130404 527474 131004 527476
rect 166404 527474 167004 527476
rect 202404 527474 203004 527476
rect 238404 527474 239004 527476
rect 274404 527474 275004 527476
rect 310404 527474 311004 527476
rect 346404 527474 347004 527476
rect 382404 527474 383004 527476
rect 418404 527474 419004 527476
rect 454404 527474 455004 527476
rect 490404 527474 491004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588080 527474 588680 527476
rect -2916 524476 -2316 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 90804 524476 91404 524478
rect 126804 524476 127404 524478
rect 162804 524476 163404 524478
rect 198804 524476 199404 524478
rect 234804 524476 235404 524478
rect 270804 524476 271404 524478
rect 306804 524476 307404 524478
rect 342804 524476 343404 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 486804 524476 487404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586240 524476 586840 524478
rect -2916 524454 586840 524476
rect -2916 524218 -2734 524454
rect -2498 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 90986 524454
rect 91222 524218 126986 524454
rect 127222 524218 162986 524454
rect 163222 524218 198986 524454
rect 199222 524218 234986 524454
rect 235222 524218 270986 524454
rect 271222 524218 306986 524454
rect 307222 524218 342986 524454
rect 343222 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586422 524454
rect 586658 524218 586840 524454
rect -2916 524134 586840 524218
rect -2916 523898 -2734 524134
rect -2498 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 90986 524134
rect 91222 523898 126986 524134
rect 127222 523898 162986 524134
rect 163222 523898 198986 524134
rect 199222 523898 234986 524134
rect 235222 523898 270986 524134
rect 271222 523898 306986 524134
rect 307222 523898 342986 524134
rect 343222 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586422 524134
rect 586658 523898 586840 524134
rect -2916 523876 586840 523898
rect -2916 523874 -2316 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 90804 523874 91404 523876
rect 126804 523874 127404 523876
rect 162804 523874 163404 523876
rect 198804 523874 199404 523876
rect 234804 523874 235404 523876
rect 270804 523874 271404 523876
rect 306804 523874 307404 523876
rect 342804 523874 343404 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 486804 523874 487404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586240 523874 586840 523876
rect -7516 517276 -6916 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 83604 517276 84204 517278
rect 119604 517276 120204 517278
rect 155604 517276 156204 517278
rect 191604 517276 192204 517278
rect 227604 517276 228204 517278
rect 263604 517276 264204 517278
rect 299604 517276 300204 517278
rect 335604 517276 336204 517278
rect 371604 517276 372204 517278
rect 407604 517276 408204 517278
rect 443604 517276 444204 517278
rect 479604 517276 480204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590840 517276 591440 517278
rect -8436 517254 592360 517276
rect -8436 517018 -7334 517254
rect -7098 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 83786 517254
rect 84022 517018 119786 517254
rect 120022 517018 155786 517254
rect 156022 517018 191786 517254
rect 192022 517018 227786 517254
rect 228022 517018 263786 517254
rect 264022 517018 299786 517254
rect 300022 517018 335786 517254
rect 336022 517018 371786 517254
rect 372022 517018 407786 517254
rect 408022 517018 443786 517254
rect 444022 517018 479786 517254
rect 480022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591022 517254
rect 591258 517018 592360 517254
rect -8436 516934 592360 517018
rect -8436 516698 -7334 516934
rect -7098 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 83786 516934
rect 84022 516698 119786 516934
rect 120022 516698 155786 516934
rect 156022 516698 191786 516934
rect 192022 516698 227786 516934
rect 228022 516698 263786 516934
rect 264022 516698 299786 516934
rect 300022 516698 335786 516934
rect 336022 516698 371786 516934
rect 372022 516698 407786 516934
rect 408022 516698 443786 516934
rect 444022 516698 479786 516934
rect 480022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591022 516934
rect 591258 516698 592360 516934
rect -8436 516676 592360 516698
rect -7516 516674 -6916 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 83604 516674 84204 516676
rect 119604 516674 120204 516676
rect 155604 516674 156204 516676
rect 191604 516674 192204 516676
rect 227604 516674 228204 516676
rect 263604 516674 264204 516676
rect 299604 516674 300204 516676
rect 335604 516674 336204 516676
rect 371604 516674 372204 516676
rect 407604 516674 408204 516676
rect 443604 516674 444204 516676
rect 479604 516674 480204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590840 516674 591440 516676
rect -5676 513676 -5076 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 80004 513676 80604 513678
rect 116004 513676 116604 513678
rect 152004 513676 152604 513678
rect 188004 513676 188604 513678
rect 224004 513676 224604 513678
rect 260004 513676 260604 513678
rect 296004 513676 296604 513678
rect 332004 513676 332604 513678
rect 368004 513676 368604 513678
rect 404004 513676 404604 513678
rect 440004 513676 440604 513678
rect 476004 513676 476604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589000 513676 589600 513678
rect -6596 513654 590520 513676
rect -6596 513418 -5494 513654
rect -5258 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 80186 513654
rect 80422 513418 116186 513654
rect 116422 513418 152186 513654
rect 152422 513418 188186 513654
rect 188422 513418 224186 513654
rect 224422 513418 260186 513654
rect 260422 513418 296186 513654
rect 296422 513418 332186 513654
rect 332422 513418 368186 513654
rect 368422 513418 404186 513654
rect 404422 513418 440186 513654
rect 440422 513418 476186 513654
rect 476422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589182 513654
rect 589418 513418 590520 513654
rect -6596 513334 590520 513418
rect -6596 513098 -5494 513334
rect -5258 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 80186 513334
rect 80422 513098 116186 513334
rect 116422 513098 152186 513334
rect 152422 513098 188186 513334
rect 188422 513098 224186 513334
rect 224422 513098 260186 513334
rect 260422 513098 296186 513334
rect 296422 513098 332186 513334
rect 332422 513098 368186 513334
rect 368422 513098 404186 513334
rect 404422 513098 440186 513334
rect 440422 513098 476186 513334
rect 476422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589182 513334
rect 589418 513098 590520 513334
rect -6596 513076 590520 513098
rect -5676 513074 -5076 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 80004 513074 80604 513076
rect 116004 513074 116604 513076
rect 152004 513074 152604 513076
rect 188004 513074 188604 513076
rect 224004 513074 224604 513076
rect 260004 513074 260604 513076
rect 296004 513074 296604 513076
rect 332004 513074 332604 513076
rect 368004 513074 368604 513076
rect 404004 513074 404604 513076
rect 440004 513074 440604 513076
rect 476004 513074 476604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589000 513074 589600 513076
rect -3836 510076 -3236 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 112404 510076 113004 510078
rect 148404 510076 149004 510078
rect 184404 510076 185004 510078
rect 220404 510076 221004 510078
rect 256404 510076 257004 510078
rect 292404 510076 293004 510078
rect 328404 510076 329004 510078
rect 364404 510076 365004 510078
rect 400404 510076 401004 510078
rect 436404 510076 437004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587160 510076 587760 510078
rect -4756 510054 588680 510076
rect -4756 509818 -3654 510054
rect -3418 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 112586 510054
rect 112822 509818 148586 510054
rect 148822 509818 184586 510054
rect 184822 509818 220586 510054
rect 220822 509818 256586 510054
rect 256822 509818 292586 510054
rect 292822 509818 328586 510054
rect 328822 509818 364586 510054
rect 364822 509818 400586 510054
rect 400822 509818 436586 510054
rect 436822 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587342 510054
rect 587578 509818 588680 510054
rect -4756 509734 588680 509818
rect -4756 509498 -3654 509734
rect -3418 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 112586 509734
rect 112822 509498 148586 509734
rect 148822 509498 184586 509734
rect 184822 509498 220586 509734
rect 220822 509498 256586 509734
rect 256822 509498 292586 509734
rect 292822 509498 328586 509734
rect 328822 509498 364586 509734
rect 364822 509498 400586 509734
rect 400822 509498 436586 509734
rect 436822 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587342 509734
rect 587578 509498 588680 509734
rect -4756 509476 588680 509498
rect -3836 509474 -3236 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 112404 509474 113004 509476
rect 148404 509474 149004 509476
rect 184404 509474 185004 509476
rect 220404 509474 221004 509476
rect 256404 509474 257004 509476
rect 292404 509474 293004 509476
rect 328404 509474 329004 509476
rect 364404 509474 365004 509476
rect 400404 509474 401004 509476
rect 436404 509474 437004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587160 509474 587760 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 108804 506476 109404 506478
rect 144804 506476 145404 506478
rect 180804 506476 181404 506478
rect 216804 506476 217404 506478
rect 252804 506476 253404 506478
rect 288804 506476 289404 506478
rect 324804 506476 325404 506478
rect 360804 506476 361404 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2916 506454 586840 506476
rect -2916 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 144986 506454
rect 145222 506218 180986 506454
rect 181222 506218 216986 506454
rect 217222 506218 252986 506454
rect 253222 506218 288986 506454
rect 289222 506218 324986 506454
rect 325222 506218 360986 506454
rect 361222 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586840 506454
rect -2916 506134 586840 506218
rect -2916 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 144986 506134
rect 145222 505898 180986 506134
rect 181222 505898 216986 506134
rect 217222 505898 252986 506134
rect 253222 505898 288986 506134
rect 289222 505898 324986 506134
rect 325222 505898 360986 506134
rect 361222 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586840 506134
rect -2916 505876 586840 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 108804 505874 109404 505876
rect 144804 505874 145404 505876
rect 180804 505874 181404 505876
rect 216804 505874 217404 505876
rect 252804 505874 253404 505876
rect 288804 505874 289404 505876
rect 324804 505874 325404 505876
rect 360804 505874 361404 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8436 499276 -7836 499278
rect 29604 499276 30204 499278
rect 65604 499276 66204 499278
rect 101604 499276 102204 499278
rect 137604 499276 138204 499278
rect 173604 499276 174204 499278
rect 209604 499276 210204 499278
rect 245604 499276 246204 499278
rect 281604 499276 282204 499278
rect 317604 499276 318204 499278
rect 353604 499276 354204 499278
rect 389604 499276 390204 499278
rect 425604 499276 426204 499278
rect 461604 499276 462204 499278
rect 497604 499276 498204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591760 499276 592360 499278
rect -8436 499254 592360 499276
rect -8436 499018 -8254 499254
rect -8018 499018 29786 499254
rect 30022 499018 65786 499254
rect 66022 499018 101786 499254
rect 102022 499018 137786 499254
rect 138022 499018 173786 499254
rect 174022 499018 209786 499254
rect 210022 499018 245786 499254
rect 246022 499018 281786 499254
rect 282022 499018 317786 499254
rect 318022 499018 353786 499254
rect 354022 499018 389786 499254
rect 390022 499018 425786 499254
rect 426022 499018 461786 499254
rect 462022 499018 497786 499254
rect 498022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 591942 499254
rect 592178 499018 592360 499254
rect -8436 498934 592360 499018
rect -8436 498698 -8254 498934
rect -8018 498698 29786 498934
rect 30022 498698 65786 498934
rect 66022 498698 101786 498934
rect 102022 498698 137786 498934
rect 138022 498698 173786 498934
rect 174022 498698 209786 498934
rect 210022 498698 245786 498934
rect 246022 498698 281786 498934
rect 282022 498698 317786 498934
rect 318022 498698 353786 498934
rect 354022 498698 389786 498934
rect 390022 498698 425786 498934
rect 426022 498698 461786 498934
rect 462022 498698 497786 498934
rect 498022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 591942 498934
rect 592178 498698 592360 498934
rect -8436 498676 592360 498698
rect -8436 498674 -7836 498676
rect 29604 498674 30204 498676
rect 65604 498674 66204 498676
rect 101604 498674 102204 498676
rect 137604 498674 138204 498676
rect 173604 498674 174204 498676
rect 209604 498674 210204 498676
rect 245604 498674 246204 498676
rect 281604 498674 282204 498676
rect 317604 498674 318204 498676
rect 353604 498674 354204 498676
rect 389604 498674 390204 498676
rect 425604 498674 426204 498676
rect 461604 498674 462204 498676
rect 497604 498674 498204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591760 498674 592360 498676
rect -6596 495676 -5996 495678
rect 26004 495676 26604 495678
rect 62004 495676 62604 495678
rect 98004 495676 98604 495678
rect 134004 495676 134604 495678
rect 170004 495676 170604 495678
rect 206004 495676 206604 495678
rect 242004 495676 242604 495678
rect 278004 495676 278604 495678
rect 314004 495676 314604 495678
rect 350004 495676 350604 495678
rect 386004 495676 386604 495678
rect 422004 495676 422604 495678
rect 458004 495676 458604 495678
rect 494004 495676 494604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 589920 495676 590520 495678
rect -6596 495654 590520 495676
rect -6596 495418 -6414 495654
rect -6178 495418 26186 495654
rect 26422 495418 62186 495654
rect 62422 495418 98186 495654
rect 98422 495418 134186 495654
rect 134422 495418 170186 495654
rect 170422 495418 206186 495654
rect 206422 495418 242186 495654
rect 242422 495418 278186 495654
rect 278422 495418 314186 495654
rect 314422 495418 350186 495654
rect 350422 495418 386186 495654
rect 386422 495418 422186 495654
rect 422422 495418 458186 495654
rect 458422 495418 494186 495654
rect 494422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590102 495654
rect 590338 495418 590520 495654
rect -6596 495334 590520 495418
rect -6596 495098 -6414 495334
rect -6178 495098 26186 495334
rect 26422 495098 62186 495334
rect 62422 495098 98186 495334
rect 98422 495098 134186 495334
rect 134422 495098 170186 495334
rect 170422 495098 206186 495334
rect 206422 495098 242186 495334
rect 242422 495098 278186 495334
rect 278422 495098 314186 495334
rect 314422 495098 350186 495334
rect 350422 495098 386186 495334
rect 386422 495098 422186 495334
rect 422422 495098 458186 495334
rect 458422 495098 494186 495334
rect 494422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590102 495334
rect 590338 495098 590520 495334
rect -6596 495076 590520 495098
rect -6596 495074 -5996 495076
rect 26004 495074 26604 495076
rect 62004 495074 62604 495076
rect 98004 495074 98604 495076
rect 134004 495074 134604 495076
rect 170004 495074 170604 495076
rect 206004 495074 206604 495076
rect 242004 495074 242604 495076
rect 278004 495074 278604 495076
rect 314004 495074 314604 495076
rect 350004 495074 350604 495076
rect 386004 495074 386604 495076
rect 422004 495074 422604 495076
rect 458004 495074 458604 495076
rect 494004 495074 494604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 589920 495074 590520 495076
rect -4756 492076 -4156 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 94404 492076 95004 492078
rect 130404 492076 131004 492078
rect 166404 492076 167004 492078
rect 202404 492076 203004 492078
rect 238404 492076 239004 492078
rect 274404 492076 275004 492078
rect 310404 492076 311004 492078
rect 346404 492076 347004 492078
rect 382404 492076 383004 492078
rect 418404 492076 419004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588080 492076 588680 492078
rect -4756 492054 588680 492076
rect -4756 491818 -4574 492054
rect -4338 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 94586 492054
rect 94822 491818 130586 492054
rect 130822 491818 166586 492054
rect 166822 491818 202586 492054
rect 202822 491818 238586 492054
rect 238822 491818 274586 492054
rect 274822 491818 310586 492054
rect 310822 491818 346586 492054
rect 346822 491818 382586 492054
rect 382822 491818 418586 492054
rect 418822 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588262 492054
rect 588498 491818 588680 492054
rect -4756 491734 588680 491818
rect -4756 491498 -4574 491734
rect -4338 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 94586 491734
rect 94822 491498 130586 491734
rect 130822 491498 166586 491734
rect 166822 491498 202586 491734
rect 202822 491498 238586 491734
rect 238822 491498 274586 491734
rect 274822 491498 310586 491734
rect 310822 491498 346586 491734
rect 346822 491498 382586 491734
rect 382822 491498 418586 491734
rect 418822 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588262 491734
rect 588498 491498 588680 491734
rect -4756 491476 588680 491498
rect -4756 491474 -4156 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 94404 491474 95004 491476
rect 130404 491474 131004 491476
rect 166404 491474 167004 491476
rect 202404 491474 203004 491476
rect 238404 491474 239004 491476
rect 274404 491474 275004 491476
rect 310404 491474 311004 491476
rect 346404 491474 347004 491476
rect 382404 491474 383004 491476
rect 418404 491474 419004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588080 491474 588680 491476
rect -2916 488476 -2316 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 162804 488476 163404 488478
rect 198804 488476 199404 488478
rect 234804 488476 235404 488478
rect 270804 488476 271404 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586240 488476 586840 488478
rect -2916 488454 586840 488476
rect -2916 488218 -2734 488454
rect -2498 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 162986 488454
rect 163222 488218 198986 488454
rect 199222 488218 234986 488454
rect 235222 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586422 488454
rect 586658 488218 586840 488454
rect -2916 488134 586840 488218
rect -2916 487898 -2734 488134
rect -2498 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 162986 488134
rect 163222 487898 198986 488134
rect 199222 487898 234986 488134
rect 235222 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586422 488134
rect 586658 487898 586840 488134
rect -2916 487876 586840 487898
rect -2916 487874 -2316 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 162804 487874 163404 487876
rect 198804 487874 199404 487876
rect 234804 487874 235404 487876
rect 270804 487874 271404 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586240 487874 586840 487876
rect -7516 481276 -6916 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 83604 481276 84204 481278
rect 119604 481276 120204 481278
rect 155604 481276 156204 481278
rect 191604 481276 192204 481278
rect 227604 481276 228204 481278
rect 263604 481276 264204 481278
rect 299604 481276 300204 481278
rect 335604 481276 336204 481278
rect 371604 481276 372204 481278
rect 407604 481276 408204 481278
rect 443604 481276 444204 481278
rect 479604 481276 480204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590840 481276 591440 481278
rect -8436 481254 592360 481276
rect -8436 481018 -7334 481254
rect -7098 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 83786 481254
rect 84022 481018 119786 481254
rect 120022 481018 155786 481254
rect 156022 481018 191786 481254
rect 192022 481018 227786 481254
rect 228022 481018 263786 481254
rect 264022 481018 299786 481254
rect 300022 481018 335786 481254
rect 336022 481018 371786 481254
rect 372022 481018 407786 481254
rect 408022 481018 443786 481254
rect 444022 481018 479786 481254
rect 480022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591022 481254
rect 591258 481018 592360 481254
rect -8436 480934 592360 481018
rect -8436 480698 -7334 480934
rect -7098 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 83786 480934
rect 84022 480698 119786 480934
rect 120022 480698 155786 480934
rect 156022 480698 191786 480934
rect 192022 480698 227786 480934
rect 228022 480698 263786 480934
rect 264022 480698 299786 480934
rect 300022 480698 335786 480934
rect 336022 480698 371786 480934
rect 372022 480698 407786 480934
rect 408022 480698 443786 480934
rect 444022 480698 479786 480934
rect 480022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591022 480934
rect 591258 480698 592360 480934
rect -8436 480676 592360 480698
rect -7516 480674 -6916 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 83604 480674 84204 480676
rect 119604 480674 120204 480676
rect 155604 480674 156204 480676
rect 191604 480674 192204 480676
rect 227604 480674 228204 480676
rect 263604 480674 264204 480676
rect 299604 480674 300204 480676
rect 335604 480674 336204 480676
rect 371604 480674 372204 480676
rect 407604 480674 408204 480676
rect 443604 480674 444204 480676
rect 479604 480674 480204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590840 480674 591440 480676
rect -5676 477676 -5076 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 80004 477676 80604 477678
rect 116004 477676 116604 477678
rect 152004 477676 152604 477678
rect 188004 477676 188604 477678
rect 224004 477676 224604 477678
rect 260004 477676 260604 477678
rect 296004 477676 296604 477678
rect 332004 477676 332604 477678
rect 368004 477676 368604 477678
rect 404004 477676 404604 477678
rect 440004 477676 440604 477678
rect 476004 477676 476604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589000 477676 589600 477678
rect -6596 477654 590520 477676
rect -6596 477418 -5494 477654
rect -5258 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 80186 477654
rect 80422 477418 116186 477654
rect 116422 477418 152186 477654
rect 152422 477418 188186 477654
rect 188422 477418 224186 477654
rect 224422 477418 260186 477654
rect 260422 477418 296186 477654
rect 296422 477418 332186 477654
rect 332422 477418 368186 477654
rect 368422 477418 404186 477654
rect 404422 477418 440186 477654
rect 440422 477418 476186 477654
rect 476422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589182 477654
rect 589418 477418 590520 477654
rect -6596 477334 590520 477418
rect -6596 477098 -5494 477334
rect -5258 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 80186 477334
rect 80422 477098 116186 477334
rect 116422 477098 152186 477334
rect 152422 477098 188186 477334
rect 188422 477098 224186 477334
rect 224422 477098 260186 477334
rect 260422 477098 296186 477334
rect 296422 477098 332186 477334
rect 332422 477098 368186 477334
rect 368422 477098 404186 477334
rect 404422 477098 440186 477334
rect 440422 477098 476186 477334
rect 476422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589182 477334
rect 589418 477098 590520 477334
rect -6596 477076 590520 477098
rect -5676 477074 -5076 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 80004 477074 80604 477076
rect 116004 477074 116604 477076
rect 152004 477074 152604 477076
rect 188004 477074 188604 477076
rect 224004 477074 224604 477076
rect 260004 477074 260604 477076
rect 296004 477074 296604 477076
rect 332004 477074 332604 477076
rect 368004 477074 368604 477076
rect 404004 477074 404604 477076
rect 440004 477074 440604 477076
rect 476004 477074 476604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589000 477074 589600 477076
rect -3836 474076 -3236 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 112404 474076 113004 474078
rect 148404 474076 149004 474078
rect 184404 474076 185004 474078
rect 220404 474076 221004 474078
rect 256404 474076 257004 474078
rect 292404 474076 293004 474078
rect 328404 474076 329004 474078
rect 364404 474076 365004 474078
rect 400404 474076 401004 474078
rect 436404 474076 437004 474078
rect 472404 474076 473004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587160 474076 587760 474078
rect -4756 474054 588680 474076
rect -4756 473818 -3654 474054
rect -3418 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 112586 474054
rect 112822 473818 148586 474054
rect 148822 473818 184586 474054
rect 184822 473818 220586 474054
rect 220822 473818 256586 474054
rect 256822 473818 292586 474054
rect 292822 473818 328586 474054
rect 328822 473818 364586 474054
rect 364822 473818 400586 474054
rect 400822 473818 436586 474054
rect 436822 473818 472586 474054
rect 472822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587342 474054
rect 587578 473818 588680 474054
rect -4756 473734 588680 473818
rect -4756 473498 -3654 473734
rect -3418 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 112586 473734
rect 112822 473498 148586 473734
rect 148822 473498 184586 473734
rect 184822 473498 220586 473734
rect 220822 473498 256586 473734
rect 256822 473498 292586 473734
rect 292822 473498 328586 473734
rect 328822 473498 364586 473734
rect 364822 473498 400586 473734
rect 400822 473498 436586 473734
rect 436822 473498 472586 473734
rect 472822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587342 473734
rect 587578 473498 588680 473734
rect -4756 473476 588680 473498
rect -3836 473474 -3236 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 112404 473474 113004 473476
rect 148404 473474 149004 473476
rect 184404 473474 185004 473476
rect 220404 473474 221004 473476
rect 256404 473474 257004 473476
rect 292404 473474 293004 473476
rect 328404 473474 329004 473476
rect 364404 473474 365004 473476
rect 400404 473474 401004 473476
rect 436404 473474 437004 473476
rect 472404 473474 473004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587160 473474 587760 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 108804 470476 109404 470478
rect 144804 470476 145404 470478
rect 180804 470476 181404 470478
rect 216804 470476 217404 470478
rect 252804 470476 253404 470478
rect 288804 470476 289404 470478
rect 324804 470476 325404 470478
rect 360804 470476 361404 470478
rect 396804 470476 397404 470478
rect 432804 470476 433404 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2916 470454 586840 470476
rect -2916 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 144986 470454
rect 145222 470218 180986 470454
rect 181222 470218 216986 470454
rect 217222 470218 252986 470454
rect 253222 470218 288986 470454
rect 289222 470218 324986 470454
rect 325222 470218 360986 470454
rect 361222 470218 396986 470454
rect 397222 470218 432986 470454
rect 433222 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586840 470454
rect -2916 470134 586840 470218
rect -2916 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 144986 470134
rect 145222 469898 180986 470134
rect 181222 469898 216986 470134
rect 217222 469898 252986 470134
rect 253222 469898 288986 470134
rect 289222 469898 324986 470134
rect 325222 469898 360986 470134
rect 361222 469898 396986 470134
rect 397222 469898 432986 470134
rect 433222 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586840 470134
rect -2916 469876 586840 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 108804 469874 109404 469876
rect 144804 469874 145404 469876
rect 180804 469874 181404 469876
rect 216804 469874 217404 469876
rect 252804 469874 253404 469876
rect 288804 469874 289404 469876
rect 324804 469874 325404 469876
rect 360804 469874 361404 469876
rect 396804 469874 397404 469876
rect 432804 469874 433404 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8436 463276 -7836 463278
rect 29604 463276 30204 463278
rect 65604 463276 66204 463278
rect 101604 463276 102204 463278
rect 137604 463276 138204 463278
rect 173604 463276 174204 463278
rect 209604 463276 210204 463278
rect 245604 463276 246204 463278
rect 281604 463276 282204 463278
rect 317604 463276 318204 463278
rect 353604 463276 354204 463278
rect 389604 463276 390204 463278
rect 425604 463276 426204 463278
rect 461604 463276 462204 463278
rect 497604 463276 498204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591760 463276 592360 463278
rect -8436 463254 592360 463276
rect -8436 463018 -8254 463254
rect -8018 463018 29786 463254
rect 30022 463018 65786 463254
rect 66022 463018 101786 463254
rect 102022 463018 137786 463254
rect 138022 463018 173786 463254
rect 174022 463018 209786 463254
rect 210022 463018 245786 463254
rect 246022 463018 281786 463254
rect 282022 463018 317786 463254
rect 318022 463018 353786 463254
rect 354022 463018 389786 463254
rect 390022 463018 425786 463254
rect 426022 463018 461786 463254
rect 462022 463018 497786 463254
rect 498022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 591942 463254
rect 592178 463018 592360 463254
rect -8436 462934 592360 463018
rect -8436 462698 -8254 462934
rect -8018 462698 29786 462934
rect 30022 462698 65786 462934
rect 66022 462698 101786 462934
rect 102022 462698 137786 462934
rect 138022 462698 173786 462934
rect 174022 462698 209786 462934
rect 210022 462698 245786 462934
rect 246022 462698 281786 462934
rect 282022 462698 317786 462934
rect 318022 462698 353786 462934
rect 354022 462698 389786 462934
rect 390022 462698 425786 462934
rect 426022 462698 461786 462934
rect 462022 462698 497786 462934
rect 498022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 591942 462934
rect 592178 462698 592360 462934
rect -8436 462676 592360 462698
rect -8436 462674 -7836 462676
rect 29604 462674 30204 462676
rect 65604 462674 66204 462676
rect 101604 462674 102204 462676
rect 137604 462674 138204 462676
rect 173604 462674 174204 462676
rect 209604 462674 210204 462676
rect 245604 462674 246204 462676
rect 281604 462674 282204 462676
rect 317604 462674 318204 462676
rect 353604 462674 354204 462676
rect 389604 462674 390204 462676
rect 425604 462674 426204 462676
rect 461604 462674 462204 462676
rect 497604 462674 498204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591760 462674 592360 462676
rect -6596 459676 -5996 459678
rect 26004 459676 26604 459678
rect 62004 459676 62604 459678
rect 98004 459676 98604 459678
rect 134004 459676 134604 459678
rect 170004 459676 170604 459678
rect 206004 459676 206604 459678
rect 242004 459676 242604 459678
rect 278004 459676 278604 459678
rect 314004 459676 314604 459678
rect 350004 459676 350604 459678
rect 386004 459676 386604 459678
rect 422004 459676 422604 459678
rect 458004 459676 458604 459678
rect 494004 459676 494604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 589920 459676 590520 459678
rect -6596 459654 590520 459676
rect -6596 459418 -6414 459654
rect -6178 459418 26186 459654
rect 26422 459418 62186 459654
rect 62422 459418 98186 459654
rect 98422 459418 134186 459654
rect 134422 459418 170186 459654
rect 170422 459418 206186 459654
rect 206422 459418 242186 459654
rect 242422 459418 278186 459654
rect 278422 459418 314186 459654
rect 314422 459418 350186 459654
rect 350422 459418 386186 459654
rect 386422 459418 422186 459654
rect 422422 459418 458186 459654
rect 458422 459418 494186 459654
rect 494422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590102 459654
rect 590338 459418 590520 459654
rect -6596 459334 590520 459418
rect -6596 459098 -6414 459334
rect -6178 459098 26186 459334
rect 26422 459098 62186 459334
rect 62422 459098 98186 459334
rect 98422 459098 134186 459334
rect 134422 459098 170186 459334
rect 170422 459098 206186 459334
rect 206422 459098 242186 459334
rect 242422 459098 278186 459334
rect 278422 459098 314186 459334
rect 314422 459098 350186 459334
rect 350422 459098 386186 459334
rect 386422 459098 422186 459334
rect 422422 459098 458186 459334
rect 458422 459098 494186 459334
rect 494422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590102 459334
rect 590338 459098 590520 459334
rect -6596 459076 590520 459098
rect -6596 459074 -5996 459076
rect 26004 459074 26604 459076
rect 62004 459074 62604 459076
rect 98004 459074 98604 459076
rect 134004 459074 134604 459076
rect 170004 459074 170604 459076
rect 206004 459074 206604 459076
rect 242004 459074 242604 459076
rect 278004 459074 278604 459076
rect 314004 459074 314604 459076
rect 350004 459074 350604 459076
rect 386004 459074 386604 459076
rect 422004 459074 422604 459076
rect 458004 459074 458604 459076
rect 494004 459074 494604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 589920 459074 590520 459076
rect -4756 456076 -4156 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 94404 456076 95004 456078
rect 130404 456076 131004 456078
rect 166404 456076 167004 456078
rect 202404 456076 203004 456078
rect 238404 456076 239004 456078
rect 274404 456076 275004 456078
rect 310404 456076 311004 456078
rect 346404 456076 347004 456078
rect 382404 456076 383004 456078
rect 418404 456076 419004 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588080 456076 588680 456078
rect -4756 456054 588680 456076
rect -4756 455818 -4574 456054
rect -4338 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 94586 456054
rect 94822 455818 130586 456054
rect 130822 455818 166586 456054
rect 166822 455818 202586 456054
rect 202822 455818 238586 456054
rect 238822 455818 274586 456054
rect 274822 455818 310586 456054
rect 310822 455818 346586 456054
rect 346822 455818 382586 456054
rect 382822 455818 418586 456054
rect 418822 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588262 456054
rect 588498 455818 588680 456054
rect -4756 455734 588680 455818
rect -4756 455498 -4574 455734
rect -4338 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 94586 455734
rect 94822 455498 130586 455734
rect 130822 455498 166586 455734
rect 166822 455498 202586 455734
rect 202822 455498 238586 455734
rect 238822 455498 274586 455734
rect 274822 455498 310586 455734
rect 310822 455498 346586 455734
rect 346822 455498 382586 455734
rect 382822 455498 418586 455734
rect 418822 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588262 455734
rect 588498 455498 588680 455734
rect -4756 455476 588680 455498
rect -4756 455474 -4156 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 94404 455474 95004 455476
rect 130404 455474 131004 455476
rect 166404 455474 167004 455476
rect 202404 455474 203004 455476
rect 238404 455474 239004 455476
rect 274404 455474 275004 455476
rect 310404 455474 311004 455476
rect 346404 455474 347004 455476
rect 382404 455474 383004 455476
rect 418404 455474 419004 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588080 455474 588680 455476
rect -2916 452476 -2316 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 162804 452476 163404 452478
rect 198804 452476 199404 452478
rect 234804 452476 235404 452478
rect 270804 452476 271404 452478
rect 306804 452476 307404 452478
rect 342804 452476 343404 452478
rect 378804 452476 379404 452478
rect 414804 452476 415404 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586240 452476 586840 452478
rect -2916 452454 586840 452476
rect -2916 452218 -2734 452454
rect -2498 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 162986 452454
rect 163222 452218 198986 452454
rect 199222 452218 234986 452454
rect 235222 452218 270986 452454
rect 271222 452218 306986 452454
rect 307222 452218 342986 452454
rect 343222 452218 378986 452454
rect 379222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586422 452454
rect 586658 452218 586840 452454
rect -2916 452134 586840 452218
rect -2916 451898 -2734 452134
rect -2498 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 162986 452134
rect 163222 451898 198986 452134
rect 199222 451898 234986 452134
rect 235222 451898 270986 452134
rect 271222 451898 306986 452134
rect 307222 451898 342986 452134
rect 343222 451898 378986 452134
rect 379222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586422 452134
rect 586658 451898 586840 452134
rect -2916 451876 586840 451898
rect -2916 451874 -2316 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 162804 451874 163404 451876
rect 198804 451874 199404 451876
rect 234804 451874 235404 451876
rect 270804 451874 271404 451876
rect 306804 451874 307404 451876
rect 342804 451874 343404 451876
rect 378804 451874 379404 451876
rect 414804 451874 415404 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586240 451874 586840 451876
rect -7516 445276 -6916 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 83604 445276 84204 445278
rect 119604 445276 120204 445278
rect 155604 445276 156204 445278
rect 191604 445276 192204 445278
rect 227604 445276 228204 445278
rect 263604 445276 264204 445278
rect 299604 445276 300204 445278
rect 335604 445276 336204 445278
rect 371604 445276 372204 445278
rect 407604 445276 408204 445278
rect 443604 445276 444204 445278
rect 479604 445276 480204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590840 445276 591440 445278
rect -8436 445254 592360 445276
rect -8436 445018 -7334 445254
rect -7098 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 83786 445254
rect 84022 445018 119786 445254
rect 120022 445018 155786 445254
rect 156022 445018 191786 445254
rect 192022 445018 227786 445254
rect 228022 445018 263786 445254
rect 264022 445018 299786 445254
rect 300022 445018 335786 445254
rect 336022 445018 371786 445254
rect 372022 445018 407786 445254
rect 408022 445018 443786 445254
rect 444022 445018 479786 445254
rect 480022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591022 445254
rect 591258 445018 592360 445254
rect -8436 444934 592360 445018
rect -8436 444698 -7334 444934
rect -7098 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 83786 444934
rect 84022 444698 119786 444934
rect 120022 444698 155786 444934
rect 156022 444698 191786 444934
rect 192022 444698 227786 444934
rect 228022 444698 263786 444934
rect 264022 444698 299786 444934
rect 300022 444698 335786 444934
rect 336022 444698 371786 444934
rect 372022 444698 407786 444934
rect 408022 444698 443786 444934
rect 444022 444698 479786 444934
rect 480022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591022 444934
rect 591258 444698 592360 444934
rect -8436 444676 592360 444698
rect -7516 444674 -6916 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 83604 444674 84204 444676
rect 119604 444674 120204 444676
rect 155604 444674 156204 444676
rect 191604 444674 192204 444676
rect 227604 444674 228204 444676
rect 263604 444674 264204 444676
rect 299604 444674 300204 444676
rect 335604 444674 336204 444676
rect 371604 444674 372204 444676
rect 407604 444674 408204 444676
rect 443604 444674 444204 444676
rect 479604 444674 480204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590840 444674 591440 444676
rect -5676 441676 -5076 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 80004 441676 80604 441678
rect 116004 441676 116604 441678
rect 152004 441676 152604 441678
rect 188004 441676 188604 441678
rect 224004 441676 224604 441678
rect 260004 441676 260604 441678
rect 296004 441676 296604 441678
rect 332004 441676 332604 441678
rect 368004 441676 368604 441678
rect 404004 441676 404604 441678
rect 440004 441676 440604 441678
rect 476004 441676 476604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589000 441676 589600 441678
rect -6596 441654 590520 441676
rect -6596 441418 -5494 441654
rect -5258 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 80186 441654
rect 80422 441418 116186 441654
rect 116422 441418 152186 441654
rect 152422 441418 188186 441654
rect 188422 441418 224186 441654
rect 224422 441418 260186 441654
rect 260422 441418 296186 441654
rect 296422 441418 332186 441654
rect 332422 441418 368186 441654
rect 368422 441418 404186 441654
rect 404422 441418 440186 441654
rect 440422 441418 476186 441654
rect 476422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589182 441654
rect 589418 441418 590520 441654
rect -6596 441334 590520 441418
rect -6596 441098 -5494 441334
rect -5258 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 80186 441334
rect 80422 441098 116186 441334
rect 116422 441098 152186 441334
rect 152422 441098 188186 441334
rect 188422 441098 224186 441334
rect 224422 441098 260186 441334
rect 260422 441098 296186 441334
rect 296422 441098 332186 441334
rect 332422 441098 368186 441334
rect 368422 441098 404186 441334
rect 404422 441098 440186 441334
rect 440422 441098 476186 441334
rect 476422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589182 441334
rect 589418 441098 590520 441334
rect -6596 441076 590520 441098
rect -5676 441074 -5076 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 80004 441074 80604 441076
rect 116004 441074 116604 441076
rect 152004 441074 152604 441076
rect 188004 441074 188604 441076
rect 224004 441074 224604 441076
rect 260004 441074 260604 441076
rect 296004 441074 296604 441076
rect 332004 441074 332604 441076
rect 368004 441074 368604 441076
rect 404004 441074 404604 441076
rect 440004 441074 440604 441076
rect 476004 441074 476604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589000 441074 589600 441076
rect -3836 438076 -3236 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 112404 438076 113004 438078
rect 148404 438076 149004 438078
rect 184404 438076 185004 438078
rect 220404 438076 221004 438078
rect 256404 438076 257004 438078
rect 292404 438076 293004 438078
rect 328404 438076 329004 438078
rect 364404 438076 365004 438078
rect 400404 438076 401004 438078
rect 436404 438076 437004 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587160 438076 587760 438078
rect -4756 438054 588680 438076
rect -4756 437818 -3654 438054
rect -3418 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 112586 438054
rect 112822 437818 148586 438054
rect 148822 437818 184586 438054
rect 184822 437818 220586 438054
rect 220822 437818 256586 438054
rect 256822 437818 292586 438054
rect 292822 437818 328586 438054
rect 328822 437818 364586 438054
rect 364822 437818 400586 438054
rect 400822 437818 436586 438054
rect 436822 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587342 438054
rect 587578 437818 588680 438054
rect -4756 437734 588680 437818
rect -4756 437498 -3654 437734
rect -3418 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 112586 437734
rect 112822 437498 148586 437734
rect 148822 437498 184586 437734
rect 184822 437498 220586 437734
rect 220822 437498 256586 437734
rect 256822 437498 292586 437734
rect 292822 437498 328586 437734
rect 328822 437498 364586 437734
rect 364822 437498 400586 437734
rect 400822 437498 436586 437734
rect 436822 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587342 437734
rect 587578 437498 588680 437734
rect -4756 437476 588680 437498
rect -3836 437474 -3236 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 112404 437474 113004 437476
rect 148404 437474 149004 437476
rect 184404 437474 185004 437476
rect 220404 437474 221004 437476
rect 256404 437474 257004 437476
rect 292404 437474 293004 437476
rect 328404 437474 329004 437476
rect 364404 437474 365004 437476
rect 400404 437474 401004 437476
rect 436404 437474 437004 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587160 437474 587760 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 108804 434476 109404 434478
rect 144804 434476 145404 434478
rect 180804 434476 181404 434478
rect 216804 434476 217404 434478
rect 252804 434476 253404 434478
rect 288804 434476 289404 434478
rect 324804 434476 325404 434478
rect 360804 434476 361404 434478
rect 396804 434476 397404 434478
rect 432804 434476 433404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2916 434454 586840 434476
rect -2916 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 144986 434454
rect 145222 434218 180986 434454
rect 181222 434218 216986 434454
rect 217222 434218 252986 434454
rect 253222 434218 288986 434454
rect 289222 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586840 434454
rect -2916 434134 586840 434218
rect -2916 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 144986 434134
rect 145222 433898 180986 434134
rect 181222 433898 216986 434134
rect 217222 433898 252986 434134
rect 253222 433898 288986 434134
rect 289222 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586840 434134
rect -2916 433876 586840 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 108804 433874 109404 433876
rect 144804 433874 145404 433876
rect 180804 433874 181404 433876
rect 216804 433874 217404 433876
rect 252804 433874 253404 433876
rect 288804 433874 289404 433876
rect 324804 433874 325404 433876
rect 360804 433874 361404 433876
rect 396804 433874 397404 433876
rect 432804 433874 433404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8436 427276 -7836 427278
rect 29604 427276 30204 427278
rect 65604 427276 66204 427278
rect 101604 427276 102204 427278
rect 137604 427276 138204 427278
rect 173604 427276 174204 427278
rect 209604 427276 210204 427278
rect 245604 427276 246204 427278
rect 281604 427276 282204 427278
rect 317604 427276 318204 427278
rect 353604 427276 354204 427278
rect 389604 427276 390204 427278
rect 425604 427276 426204 427278
rect 461604 427276 462204 427278
rect 497604 427276 498204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591760 427276 592360 427278
rect -8436 427254 592360 427276
rect -8436 427018 -8254 427254
rect -8018 427018 29786 427254
rect 30022 427018 65786 427254
rect 66022 427018 101786 427254
rect 102022 427018 137786 427254
rect 138022 427018 173786 427254
rect 174022 427018 209786 427254
rect 210022 427018 245786 427254
rect 246022 427018 281786 427254
rect 282022 427018 317786 427254
rect 318022 427018 353786 427254
rect 354022 427018 389786 427254
rect 390022 427018 425786 427254
rect 426022 427018 461786 427254
rect 462022 427018 497786 427254
rect 498022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 591942 427254
rect 592178 427018 592360 427254
rect -8436 426934 592360 427018
rect -8436 426698 -8254 426934
rect -8018 426698 29786 426934
rect 30022 426698 65786 426934
rect 66022 426698 101786 426934
rect 102022 426698 137786 426934
rect 138022 426698 173786 426934
rect 174022 426698 209786 426934
rect 210022 426698 245786 426934
rect 246022 426698 281786 426934
rect 282022 426698 317786 426934
rect 318022 426698 353786 426934
rect 354022 426698 389786 426934
rect 390022 426698 425786 426934
rect 426022 426698 461786 426934
rect 462022 426698 497786 426934
rect 498022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 591942 426934
rect 592178 426698 592360 426934
rect -8436 426676 592360 426698
rect -8436 426674 -7836 426676
rect 29604 426674 30204 426676
rect 65604 426674 66204 426676
rect 101604 426674 102204 426676
rect 137604 426674 138204 426676
rect 173604 426674 174204 426676
rect 209604 426674 210204 426676
rect 245604 426674 246204 426676
rect 281604 426674 282204 426676
rect 317604 426674 318204 426676
rect 353604 426674 354204 426676
rect 389604 426674 390204 426676
rect 425604 426674 426204 426676
rect 461604 426674 462204 426676
rect 497604 426674 498204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591760 426674 592360 426676
rect -6596 423676 -5996 423678
rect 26004 423676 26604 423678
rect 62004 423676 62604 423678
rect 98004 423676 98604 423678
rect 134004 423676 134604 423678
rect 170004 423676 170604 423678
rect 206004 423676 206604 423678
rect 242004 423676 242604 423678
rect 278004 423676 278604 423678
rect 314004 423676 314604 423678
rect 350004 423676 350604 423678
rect 386004 423676 386604 423678
rect 422004 423676 422604 423678
rect 458004 423676 458604 423678
rect 494004 423676 494604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 589920 423676 590520 423678
rect -6596 423654 590520 423676
rect -6596 423418 -6414 423654
rect -6178 423418 26186 423654
rect 26422 423418 62186 423654
rect 62422 423418 98186 423654
rect 98422 423418 134186 423654
rect 134422 423418 170186 423654
rect 170422 423418 206186 423654
rect 206422 423418 242186 423654
rect 242422 423418 278186 423654
rect 278422 423418 314186 423654
rect 314422 423418 350186 423654
rect 350422 423418 386186 423654
rect 386422 423418 422186 423654
rect 422422 423418 458186 423654
rect 458422 423418 494186 423654
rect 494422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590102 423654
rect 590338 423418 590520 423654
rect -6596 423334 590520 423418
rect -6596 423098 -6414 423334
rect -6178 423098 26186 423334
rect 26422 423098 62186 423334
rect 62422 423098 98186 423334
rect 98422 423098 134186 423334
rect 134422 423098 170186 423334
rect 170422 423098 206186 423334
rect 206422 423098 242186 423334
rect 242422 423098 278186 423334
rect 278422 423098 314186 423334
rect 314422 423098 350186 423334
rect 350422 423098 386186 423334
rect 386422 423098 422186 423334
rect 422422 423098 458186 423334
rect 458422 423098 494186 423334
rect 494422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590102 423334
rect 590338 423098 590520 423334
rect -6596 423076 590520 423098
rect -6596 423074 -5996 423076
rect 26004 423074 26604 423076
rect 62004 423074 62604 423076
rect 98004 423074 98604 423076
rect 134004 423074 134604 423076
rect 170004 423074 170604 423076
rect 206004 423074 206604 423076
rect 242004 423074 242604 423076
rect 278004 423074 278604 423076
rect 314004 423074 314604 423076
rect 350004 423074 350604 423076
rect 386004 423074 386604 423076
rect 422004 423074 422604 423076
rect 458004 423074 458604 423076
rect 494004 423074 494604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 589920 423074 590520 423076
rect -4756 420076 -4156 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 94404 420076 95004 420078
rect 130404 420076 131004 420078
rect 166404 420076 167004 420078
rect 202404 420076 203004 420078
rect 238404 420076 239004 420078
rect 274404 420076 275004 420078
rect 310404 420076 311004 420078
rect 346404 420076 347004 420078
rect 382404 420076 383004 420078
rect 418404 420076 419004 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588080 420076 588680 420078
rect -4756 420054 588680 420076
rect -4756 419818 -4574 420054
rect -4338 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 94586 420054
rect 94822 419818 130586 420054
rect 130822 419818 166586 420054
rect 166822 419818 202586 420054
rect 202822 419818 238586 420054
rect 238822 419818 274586 420054
rect 274822 419818 310586 420054
rect 310822 419818 346586 420054
rect 346822 419818 382586 420054
rect 382822 419818 418586 420054
rect 418822 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588262 420054
rect 588498 419818 588680 420054
rect -4756 419734 588680 419818
rect -4756 419498 -4574 419734
rect -4338 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 94586 419734
rect 94822 419498 130586 419734
rect 130822 419498 166586 419734
rect 166822 419498 202586 419734
rect 202822 419498 238586 419734
rect 238822 419498 274586 419734
rect 274822 419498 310586 419734
rect 310822 419498 346586 419734
rect 346822 419498 382586 419734
rect 382822 419498 418586 419734
rect 418822 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588262 419734
rect 588498 419498 588680 419734
rect -4756 419476 588680 419498
rect -4756 419474 -4156 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 94404 419474 95004 419476
rect 130404 419474 131004 419476
rect 166404 419474 167004 419476
rect 202404 419474 203004 419476
rect 238404 419474 239004 419476
rect 274404 419474 275004 419476
rect 310404 419474 311004 419476
rect 346404 419474 347004 419476
rect 382404 419474 383004 419476
rect 418404 419474 419004 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588080 419474 588680 419476
rect -2916 416476 -2316 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 90804 416476 91404 416478
rect 126804 416476 127404 416478
rect 162804 416476 163404 416478
rect 198804 416476 199404 416478
rect 234804 416476 235404 416478
rect 270804 416476 271404 416478
rect 306804 416476 307404 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586240 416476 586840 416478
rect -2916 416454 586840 416476
rect -2916 416218 -2734 416454
rect -2498 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 90986 416454
rect 91222 416218 126986 416454
rect 127222 416218 162986 416454
rect 163222 416218 198986 416454
rect 199222 416218 234986 416454
rect 235222 416218 270986 416454
rect 271222 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586422 416454
rect 586658 416218 586840 416454
rect -2916 416134 586840 416218
rect -2916 415898 -2734 416134
rect -2498 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 90986 416134
rect 91222 415898 126986 416134
rect 127222 415898 162986 416134
rect 163222 415898 198986 416134
rect 199222 415898 234986 416134
rect 235222 415898 270986 416134
rect 271222 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586422 416134
rect 586658 415898 586840 416134
rect -2916 415876 586840 415898
rect -2916 415874 -2316 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 90804 415874 91404 415876
rect 126804 415874 127404 415876
rect 162804 415874 163404 415876
rect 198804 415874 199404 415876
rect 234804 415874 235404 415876
rect 270804 415874 271404 415876
rect 306804 415874 307404 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586240 415874 586840 415876
rect -7516 409276 -6916 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 83604 409276 84204 409278
rect 119604 409276 120204 409278
rect 155604 409276 156204 409278
rect 191604 409276 192204 409278
rect 227604 409276 228204 409278
rect 263604 409276 264204 409278
rect 299604 409276 300204 409278
rect 335604 409276 336204 409278
rect 371604 409276 372204 409278
rect 407604 409276 408204 409278
rect 443604 409276 444204 409278
rect 479604 409276 480204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590840 409276 591440 409278
rect -8436 409254 592360 409276
rect -8436 409018 -7334 409254
rect -7098 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 83786 409254
rect 84022 409018 119786 409254
rect 120022 409018 155786 409254
rect 156022 409018 191786 409254
rect 192022 409018 227786 409254
rect 228022 409018 263786 409254
rect 264022 409018 299786 409254
rect 300022 409018 335786 409254
rect 336022 409018 371786 409254
rect 372022 409018 407786 409254
rect 408022 409018 443786 409254
rect 444022 409018 479786 409254
rect 480022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591022 409254
rect 591258 409018 592360 409254
rect -8436 408934 592360 409018
rect -8436 408698 -7334 408934
rect -7098 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 83786 408934
rect 84022 408698 119786 408934
rect 120022 408698 155786 408934
rect 156022 408698 191786 408934
rect 192022 408698 227786 408934
rect 228022 408698 263786 408934
rect 264022 408698 299786 408934
rect 300022 408698 335786 408934
rect 336022 408698 371786 408934
rect 372022 408698 407786 408934
rect 408022 408698 443786 408934
rect 444022 408698 479786 408934
rect 480022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591022 408934
rect 591258 408698 592360 408934
rect -8436 408676 592360 408698
rect -7516 408674 -6916 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 83604 408674 84204 408676
rect 119604 408674 120204 408676
rect 155604 408674 156204 408676
rect 191604 408674 192204 408676
rect 227604 408674 228204 408676
rect 263604 408674 264204 408676
rect 299604 408674 300204 408676
rect 335604 408674 336204 408676
rect 371604 408674 372204 408676
rect 407604 408674 408204 408676
rect 443604 408674 444204 408676
rect 479604 408674 480204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590840 408674 591440 408676
rect -5676 405676 -5076 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 80004 405676 80604 405678
rect 116004 405676 116604 405678
rect 152004 405676 152604 405678
rect 188004 405676 188604 405678
rect 224004 405676 224604 405678
rect 260004 405676 260604 405678
rect 296004 405676 296604 405678
rect 332004 405676 332604 405678
rect 368004 405676 368604 405678
rect 404004 405676 404604 405678
rect 440004 405676 440604 405678
rect 476004 405676 476604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589000 405676 589600 405678
rect -6596 405654 590520 405676
rect -6596 405418 -5494 405654
rect -5258 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 80186 405654
rect 80422 405418 116186 405654
rect 116422 405418 152186 405654
rect 152422 405418 188186 405654
rect 188422 405418 224186 405654
rect 224422 405418 260186 405654
rect 260422 405418 296186 405654
rect 296422 405418 332186 405654
rect 332422 405418 368186 405654
rect 368422 405418 404186 405654
rect 404422 405418 440186 405654
rect 440422 405418 476186 405654
rect 476422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589182 405654
rect 589418 405418 590520 405654
rect -6596 405334 590520 405418
rect -6596 405098 -5494 405334
rect -5258 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 80186 405334
rect 80422 405098 116186 405334
rect 116422 405098 152186 405334
rect 152422 405098 188186 405334
rect 188422 405098 224186 405334
rect 224422 405098 260186 405334
rect 260422 405098 296186 405334
rect 296422 405098 332186 405334
rect 332422 405098 368186 405334
rect 368422 405098 404186 405334
rect 404422 405098 440186 405334
rect 440422 405098 476186 405334
rect 476422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589182 405334
rect 589418 405098 590520 405334
rect -6596 405076 590520 405098
rect -5676 405074 -5076 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 80004 405074 80604 405076
rect 116004 405074 116604 405076
rect 152004 405074 152604 405076
rect 188004 405074 188604 405076
rect 224004 405074 224604 405076
rect 260004 405074 260604 405076
rect 296004 405074 296604 405076
rect 332004 405074 332604 405076
rect 368004 405074 368604 405076
rect 404004 405074 404604 405076
rect 440004 405074 440604 405076
rect 476004 405074 476604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589000 405074 589600 405076
rect -3836 402076 -3236 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 112404 402076 113004 402078
rect 148404 402076 149004 402078
rect 184404 402076 185004 402078
rect 220404 402076 221004 402078
rect 256404 402076 257004 402078
rect 292404 402076 293004 402078
rect 328404 402076 329004 402078
rect 364404 402076 365004 402078
rect 400404 402076 401004 402078
rect 436404 402076 437004 402078
rect 472404 402076 473004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587160 402076 587760 402078
rect -4756 402054 588680 402076
rect -4756 401818 -3654 402054
rect -3418 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 112586 402054
rect 112822 401818 148586 402054
rect 148822 401818 184586 402054
rect 184822 401818 220586 402054
rect 220822 401818 256586 402054
rect 256822 401818 292586 402054
rect 292822 401818 328586 402054
rect 328822 401818 364586 402054
rect 364822 401818 400586 402054
rect 400822 401818 436586 402054
rect 436822 401818 472586 402054
rect 472822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587342 402054
rect 587578 401818 588680 402054
rect -4756 401734 588680 401818
rect -4756 401498 -3654 401734
rect -3418 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 112586 401734
rect 112822 401498 148586 401734
rect 148822 401498 184586 401734
rect 184822 401498 220586 401734
rect 220822 401498 256586 401734
rect 256822 401498 292586 401734
rect 292822 401498 328586 401734
rect 328822 401498 364586 401734
rect 364822 401498 400586 401734
rect 400822 401498 436586 401734
rect 436822 401498 472586 401734
rect 472822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587342 401734
rect 587578 401498 588680 401734
rect -4756 401476 588680 401498
rect -3836 401474 -3236 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 112404 401474 113004 401476
rect 148404 401474 149004 401476
rect 184404 401474 185004 401476
rect 220404 401474 221004 401476
rect 256404 401474 257004 401476
rect 292404 401474 293004 401476
rect 328404 401474 329004 401476
rect 364404 401474 365004 401476
rect 400404 401474 401004 401476
rect 436404 401474 437004 401476
rect 472404 401474 473004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587160 401474 587760 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 144804 398476 145404 398478
rect 180804 398476 181404 398478
rect 216804 398476 217404 398478
rect 252804 398476 253404 398478
rect 288804 398476 289404 398478
rect 324804 398476 325404 398478
rect 360804 398476 361404 398478
rect 396804 398476 397404 398478
rect 432804 398476 433404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2916 398454 586840 398476
rect -2916 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 144986 398454
rect 145222 398218 180986 398454
rect 181222 398218 216986 398454
rect 217222 398218 252986 398454
rect 253222 398218 288986 398454
rect 289222 398218 324986 398454
rect 325222 398218 360986 398454
rect 361222 398218 396986 398454
rect 397222 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586840 398454
rect -2916 398134 586840 398218
rect -2916 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 144986 398134
rect 145222 397898 180986 398134
rect 181222 397898 216986 398134
rect 217222 397898 252986 398134
rect 253222 397898 288986 398134
rect 289222 397898 324986 398134
rect 325222 397898 360986 398134
rect 361222 397898 396986 398134
rect 397222 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586840 398134
rect -2916 397876 586840 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 144804 397874 145404 397876
rect 180804 397874 181404 397876
rect 216804 397874 217404 397876
rect 252804 397874 253404 397876
rect 288804 397874 289404 397876
rect 324804 397874 325404 397876
rect 360804 397874 361404 397876
rect 396804 397874 397404 397876
rect 432804 397874 433404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8436 391276 -7836 391278
rect 29604 391276 30204 391278
rect 65604 391276 66204 391278
rect 101604 391276 102204 391278
rect 137604 391276 138204 391278
rect 173604 391276 174204 391278
rect 209604 391276 210204 391278
rect 245604 391276 246204 391278
rect 281604 391276 282204 391278
rect 317604 391276 318204 391278
rect 353604 391276 354204 391278
rect 389604 391276 390204 391278
rect 425604 391276 426204 391278
rect 461604 391276 462204 391278
rect 497604 391276 498204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591760 391276 592360 391278
rect -8436 391254 592360 391276
rect -8436 391018 -8254 391254
rect -8018 391018 29786 391254
rect 30022 391018 65786 391254
rect 66022 391018 101786 391254
rect 102022 391018 137786 391254
rect 138022 391018 173786 391254
rect 174022 391018 209786 391254
rect 210022 391018 245786 391254
rect 246022 391018 281786 391254
rect 282022 391018 317786 391254
rect 318022 391018 353786 391254
rect 354022 391018 389786 391254
rect 390022 391018 425786 391254
rect 426022 391018 461786 391254
rect 462022 391018 497786 391254
rect 498022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 591942 391254
rect 592178 391018 592360 391254
rect -8436 390934 592360 391018
rect -8436 390698 -8254 390934
rect -8018 390698 29786 390934
rect 30022 390698 65786 390934
rect 66022 390698 101786 390934
rect 102022 390698 137786 390934
rect 138022 390698 173786 390934
rect 174022 390698 209786 390934
rect 210022 390698 245786 390934
rect 246022 390698 281786 390934
rect 282022 390698 317786 390934
rect 318022 390698 353786 390934
rect 354022 390698 389786 390934
rect 390022 390698 425786 390934
rect 426022 390698 461786 390934
rect 462022 390698 497786 390934
rect 498022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 591942 390934
rect 592178 390698 592360 390934
rect -8436 390676 592360 390698
rect -8436 390674 -7836 390676
rect 29604 390674 30204 390676
rect 65604 390674 66204 390676
rect 101604 390674 102204 390676
rect 137604 390674 138204 390676
rect 173604 390674 174204 390676
rect 209604 390674 210204 390676
rect 245604 390674 246204 390676
rect 281604 390674 282204 390676
rect 317604 390674 318204 390676
rect 353604 390674 354204 390676
rect 389604 390674 390204 390676
rect 425604 390674 426204 390676
rect 461604 390674 462204 390676
rect 497604 390674 498204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591760 390674 592360 390676
rect -6596 387676 -5996 387678
rect 26004 387676 26604 387678
rect 62004 387676 62604 387678
rect 98004 387676 98604 387678
rect 134004 387676 134604 387678
rect 170004 387676 170604 387678
rect 206004 387676 206604 387678
rect 242004 387676 242604 387678
rect 278004 387676 278604 387678
rect 314004 387676 314604 387678
rect 350004 387676 350604 387678
rect 386004 387676 386604 387678
rect 422004 387676 422604 387678
rect 458004 387676 458604 387678
rect 494004 387676 494604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 589920 387676 590520 387678
rect -6596 387654 590520 387676
rect -6596 387418 -6414 387654
rect -6178 387418 26186 387654
rect 26422 387418 62186 387654
rect 62422 387418 98186 387654
rect 98422 387418 134186 387654
rect 134422 387418 170186 387654
rect 170422 387418 206186 387654
rect 206422 387418 242186 387654
rect 242422 387418 278186 387654
rect 278422 387418 314186 387654
rect 314422 387418 350186 387654
rect 350422 387418 386186 387654
rect 386422 387418 422186 387654
rect 422422 387418 458186 387654
rect 458422 387418 494186 387654
rect 494422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590102 387654
rect 590338 387418 590520 387654
rect -6596 387334 590520 387418
rect -6596 387098 -6414 387334
rect -6178 387098 26186 387334
rect 26422 387098 62186 387334
rect 62422 387098 98186 387334
rect 98422 387098 134186 387334
rect 134422 387098 170186 387334
rect 170422 387098 206186 387334
rect 206422 387098 242186 387334
rect 242422 387098 278186 387334
rect 278422 387098 314186 387334
rect 314422 387098 350186 387334
rect 350422 387098 386186 387334
rect 386422 387098 422186 387334
rect 422422 387098 458186 387334
rect 458422 387098 494186 387334
rect 494422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590102 387334
rect 590338 387098 590520 387334
rect -6596 387076 590520 387098
rect -6596 387074 -5996 387076
rect 26004 387074 26604 387076
rect 62004 387074 62604 387076
rect 98004 387074 98604 387076
rect 134004 387074 134604 387076
rect 170004 387074 170604 387076
rect 206004 387074 206604 387076
rect 242004 387074 242604 387076
rect 278004 387074 278604 387076
rect 314004 387074 314604 387076
rect 350004 387074 350604 387076
rect 386004 387074 386604 387076
rect 422004 387074 422604 387076
rect 458004 387074 458604 387076
rect 494004 387074 494604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 589920 387074 590520 387076
rect -4756 384076 -4156 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 94404 384076 95004 384078
rect 130404 384076 131004 384078
rect 166404 384076 167004 384078
rect 202404 384076 203004 384078
rect 238404 384076 239004 384078
rect 274404 384076 275004 384078
rect 310404 384076 311004 384078
rect 346404 384076 347004 384078
rect 382404 384076 383004 384078
rect 418404 384076 419004 384078
rect 454404 384076 455004 384078
rect 490404 384076 491004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588080 384076 588680 384078
rect -4756 384054 588680 384076
rect -4756 383818 -4574 384054
rect -4338 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 94586 384054
rect 94822 383818 130586 384054
rect 130822 383818 166586 384054
rect 166822 383818 202586 384054
rect 202822 383818 238586 384054
rect 238822 383818 274586 384054
rect 274822 383818 310586 384054
rect 310822 383818 346586 384054
rect 346822 383818 382586 384054
rect 382822 383818 418586 384054
rect 418822 383818 454586 384054
rect 454822 383818 490586 384054
rect 490822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588262 384054
rect 588498 383818 588680 384054
rect -4756 383734 588680 383818
rect -4756 383498 -4574 383734
rect -4338 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 94586 383734
rect 94822 383498 130586 383734
rect 130822 383498 166586 383734
rect 166822 383498 202586 383734
rect 202822 383498 238586 383734
rect 238822 383498 274586 383734
rect 274822 383498 310586 383734
rect 310822 383498 346586 383734
rect 346822 383498 382586 383734
rect 382822 383498 418586 383734
rect 418822 383498 454586 383734
rect 454822 383498 490586 383734
rect 490822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588262 383734
rect 588498 383498 588680 383734
rect -4756 383476 588680 383498
rect -4756 383474 -4156 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 94404 383474 95004 383476
rect 130404 383474 131004 383476
rect 166404 383474 167004 383476
rect 202404 383474 203004 383476
rect 238404 383474 239004 383476
rect 274404 383474 275004 383476
rect 310404 383474 311004 383476
rect 346404 383474 347004 383476
rect 382404 383474 383004 383476
rect 418404 383474 419004 383476
rect 454404 383474 455004 383476
rect 490404 383474 491004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588080 383474 588680 383476
rect -2916 380476 -2316 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 162804 380476 163404 380478
rect 198804 380476 199404 380478
rect 234804 380476 235404 380478
rect 270804 380476 271404 380478
rect 306804 380476 307404 380478
rect 342804 380476 343404 380478
rect 378804 380476 379404 380478
rect 414804 380476 415404 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586240 380476 586840 380478
rect -2916 380454 586840 380476
rect -2916 380218 -2734 380454
rect -2498 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 198986 380454
rect 199222 380218 234986 380454
rect 235222 380218 270986 380454
rect 271222 380218 306986 380454
rect 307222 380218 342986 380454
rect 343222 380218 378986 380454
rect 379222 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586422 380454
rect 586658 380218 586840 380454
rect -2916 380134 586840 380218
rect -2916 379898 -2734 380134
rect -2498 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 198986 380134
rect 199222 379898 234986 380134
rect 235222 379898 270986 380134
rect 271222 379898 306986 380134
rect 307222 379898 342986 380134
rect 343222 379898 378986 380134
rect 379222 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586422 380134
rect 586658 379898 586840 380134
rect -2916 379876 586840 379898
rect -2916 379874 -2316 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 162804 379874 163404 379876
rect 198804 379874 199404 379876
rect 234804 379874 235404 379876
rect 270804 379874 271404 379876
rect 306804 379874 307404 379876
rect 342804 379874 343404 379876
rect 378804 379874 379404 379876
rect 414804 379874 415404 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586240 379874 586840 379876
rect -7516 373276 -6916 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 83604 373276 84204 373278
rect 119604 373276 120204 373278
rect 155604 373276 156204 373278
rect 191604 373276 192204 373278
rect 227604 373276 228204 373278
rect 263604 373276 264204 373278
rect 299604 373276 300204 373278
rect 335604 373276 336204 373278
rect 371604 373276 372204 373278
rect 407604 373276 408204 373278
rect 443604 373276 444204 373278
rect 479604 373276 480204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590840 373276 591440 373278
rect -8436 373254 592360 373276
rect -8436 373018 -7334 373254
rect -7098 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 83786 373254
rect 84022 373018 119786 373254
rect 120022 373018 155786 373254
rect 156022 373018 191786 373254
rect 192022 373018 227786 373254
rect 228022 373018 263786 373254
rect 264022 373018 299786 373254
rect 300022 373018 335786 373254
rect 336022 373018 371786 373254
rect 372022 373018 407786 373254
rect 408022 373018 443786 373254
rect 444022 373018 479786 373254
rect 480022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591022 373254
rect 591258 373018 592360 373254
rect -8436 372934 592360 373018
rect -8436 372698 -7334 372934
rect -7098 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 83786 372934
rect 84022 372698 119786 372934
rect 120022 372698 155786 372934
rect 156022 372698 191786 372934
rect 192022 372698 227786 372934
rect 228022 372698 263786 372934
rect 264022 372698 299786 372934
rect 300022 372698 335786 372934
rect 336022 372698 371786 372934
rect 372022 372698 407786 372934
rect 408022 372698 443786 372934
rect 444022 372698 479786 372934
rect 480022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591022 372934
rect 591258 372698 592360 372934
rect -8436 372676 592360 372698
rect -7516 372674 -6916 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 83604 372674 84204 372676
rect 119604 372674 120204 372676
rect 155604 372674 156204 372676
rect 191604 372674 192204 372676
rect 227604 372674 228204 372676
rect 263604 372674 264204 372676
rect 299604 372674 300204 372676
rect 335604 372674 336204 372676
rect 371604 372674 372204 372676
rect 407604 372674 408204 372676
rect 443604 372674 444204 372676
rect 479604 372674 480204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590840 372674 591440 372676
rect -5676 369676 -5076 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 80004 369676 80604 369678
rect 116004 369676 116604 369678
rect 152004 369676 152604 369678
rect 188004 369676 188604 369678
rect 224004 369676 224604 369678
rect 260004 369676 260604 369678
rect 296004 369676 296604 369678
rect 332004 369676 332604 369678
rect 368004 369676 368604 369678
rect 404004 369676 404604 369678
rect 440004 369676 440604 369678
rect 476004 369676 476604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589000 369676 589600 369678
rect -6596 369654 590520 369676
rect -6596 369418 -5494 369654
rect -5258 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 80186 369654
rect 80422 369418 116186 369654
rect 116422 369418 152186 369654
rect 152422 369418 188186 369654
rect 188422 369418 224186 369654
rect 224422 369418 260186 369654
rect 260422 369418 296186 369654
rect 296422 369418 332186 369654
rect 332422 369418 368186 369654
rect 368422 369418 404186 369654
rect 404422 369418 440186 369654
rect 440422 369418 476186 369654
rect 476422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589182 369654
rect 589418 369418 590520 369654
rect -6596 369334 590520 369418
rect -6596 369098 -5494 369334
rect -5258 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 80186 369334
rect 80422 369098 116186 369334
rect 116422 369098 152186 369334
rect 152422 369098 188186 369334
rect 188422 369098 224186 369334
rect 224422 369098 260186 369334
rect 260422 369098 296186 369334
rect 296422 369098 332186 369334
rect 332422 369098 368186 369334
rect 368422 369098 404186 369334
rect 404422 369098 440186 369334
rect 440422 369098 476186 369334
rect 476422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589182 369334
rect 589418 369098 590520 369334
rect -6596 369076 590520 369098
rect -5676 369074 -5076 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 80004 369074 80604 369076
rect 116004 369074 116604 369076
rect 152004 369074 152604 369076
rect 188004 369074 188604 369076
rect 224004 369074 224604 369076
rect 260004 369074 260604 369076
rect 296004 369074 296604 369076
rect 332004 369074 332604 369076
rect 368004 369074 368604 369076
rect 404004 369074 404604 369076
rect 440004 369074 440604 369076
rect 476004 369074 476604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589000 369074 589600 369076
rect -3836 366076 -3236 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 76404 366076 77004 366078
rect 112404 366076 113004 366078
rect 148404 366076 149004 366078
rect 184404 366076 185004 366078
rect 220404 366076 221004 366078
rect 256404 366076 257004 366078
rect 292404 366076 293004 366078
rect 328404 366076 329004 366078
rect 364404 366076 365004 366078
rect 400404 366076 401004 366078
rect 436404 366076 437004 366078
rect 472404 366076 473004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587160 366076 587760 366078
rect -4756 366054 588680 366076
rect -4756 365818 -3654 366054
rect -3418 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 76586 366054
rect 76822 365818 112586 366054
rect 112822 365818 148586 366054
rect 148822 365818 184586 366054
rect 184822 365818 220586 366054
rect 220822 365818 256586 366054
rect 256822 365818 292586 366054
rect 292822 365818 328586 366054
rect 328822 365818 364586 366054
rect 364822 365818 400586 366054
rect 400822 365818 436586 366054
rect 436822 365818 472586 366054
rect 472822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587342 366054
rect 587578 365818 588680 366054
rect -4756 365734 588680 365818
rect -4756 365498 -3654 365734
rect -3418 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 76586 365734
rect 76822 365498 112586 365734
rect 112822 365498 148586 365734
rect 148822 365498 184586 365734
rect 184822 365498 220586 365734
rect 220822 365498 256586 365734
rect 256822 365498 292586 365734
rect 292822 365498 328586 365734
rect 328822 365498 364586 365734
rect 364822 365498 400586 365734
rect 400822 365498 436586 365734
rect 436822 365498 472586 365734
rect 472822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587342 365734
rect 587578 365498 588680 365734
rect -4756 365476 588680 365498
rect -3836 365474 -3236 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 76404 365474 77004 365476
rect 112404 365474 113004 365476
rect 148404 365474 149004 365476
rect 184404 365474 185004 365476
rect 220404 365474 221004 365476
rect 256404 365474 257004 365476
rect 292404 365474 293004 365476
rect 328404 365474 329004 365476
rect 364404 365474 365004 365476
rect 400404 365474 401004 365476
rect 436404 365474 437004 365476
rect 472404 365474 473004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587160 365474 587760 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 108804 362476 109404 362478
rect 144804 362476 145404 362478
rect 180804 362476 181404 362478
rect 216804 362476 217404 362478
rect 252804 362476 253404 362478
rect 288804 362476 289404 362478
rect 324804 362476 325404 362478
rect 360804 362476 361404 362478
rect 396804 362476 397404 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2916 362454 586840 362476
rect -2916 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 216986 362454
rect 217222 362218 252986 362454
rect 253222 362218 288986 362454
rect 289222 362218 324986 362454
rect 325222 362218 360986 362454
rect 361222 362218 396986 362454
rect 397222 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586840 362454
rect -2916 362134 586840 362218
rect -2916 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 216986 362134
rect 217222 361898 252986 362134
rect 253222 361898 288986 362134
rect 289222 361898 324986 362134
rect 325222 361898 360986 362134
rect 361222 361898 396986 362134
rect 397222 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586840 362134
rect -2916 361876 586840 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 108804 361874 109404 361876
rect 144804 361874 145404 361876
rect 180804 361874 181404 361876
rect 216804 361874 217404 361876
rect 252804 361874 253404 361876
rect 288804 361874 289404 361876
rect 324804 361874 325404 361876
rect 360804 361874 361404 361876
rect 396804 361874 397404 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8436 355276 -7836 355278
rect 29604 355276 30204 355278
rect 65604 355276 66204 355278
rect 101604 355276 102204 355278
rect 137604 355276 138204 355278
rect 173604 355276 174204 355278
rect 209604 355276 210204 355278
rect 245604 355276 246204 355278
rect 281604 355276 282204 355278
rect 317604 355276 318204 355278
rect 353604 355276 354204 355278
rect 389604 355276 390204 355278
rect 425604 355276 426204 355278
rect 461604 355276 462204 355278
rect 497604 355276 498204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591760 355276 592360 355278
rect -8436 355254 592360 355276
rect -8436 355018 -8254 355254
rect -8018 355018 29786 355254
rect 30022 355018 65786 355254
rect 66022 355018 101786 355254
rect 102022 355018 137786 355254
rect 138022 355018 173786 355254
rect 174022 355018 209786 355254
rect 210022 355018 245786 355254
rect 246022 355018 281786 355254
rect 282022 355018 317786 355254
rect 318022 355018 353786 355254
rect 354022 355018 389786 355254
rect 390022 355018 425786 355254
rect 426022 355018 461786 355254
rect 462022 355018 497786 355254
rect 498022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 591942 355254
rect 592178 355018 592360 355254
rect -8436 354934 592360 355018
rect -8436 354698 -8254 354934
rect -8018 354698 29786 354934
rect 30022 354698 65786 354934
rect 66022 354698 101786 354934
rect 102022 354698 137786 354934
rect 138022 354698 173786 354934
rect 174022 354698 209786 354934
rect 210022 354698 245786 354934
rect 246022 354698 281786 354934
rect 282022 354698 317786 354934
rect 318022 354698 353786 354934
rect 354022 354698 389786 354934
rect 390022 354698 425786 354934
rect 426022 354698 461786 354934
rect 462022 354698 497786 354934
rect 498022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 591942 354934
rect 592178 354698 592360 354934
rect -8436 354676 592360 354698
rect -8436 354674 -7836 354676
rect 29604 354674 30204 354676
rect 65604 354674 66204 354676
rect 101604 354674 102204 354676
rect 137604 354674 138204 354676
rect 173604 354674 174204 354676
rect 209604 354674 210204 354676
rect 245604 354674 246204 354676
rect 281604 354674 282204 354676
rect 317604 354674 318204 354676
rect 353604 354674 354204 354676
rect 389604 354674 390204 354676
rect 425604 354674 426204 354676
rect 461604 354674 462204 354676
rect 497604 354674 498204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591760 354674 592360 354676
rect -6596 351676 -5996 351678
rect 26004 351676 26604 351678
rect 62004 351676 62604 351678
rect 98004 351676 98604 351678
rect 134004 351676 134604 351678
rect 170004 351676 170604 351678
rect 206004 351676 206604 351678
rect 242004 351676 242604 351678
rect 278004 351676 278604 351678
rect 314004 351676 314604 351678
rect 350004 351676 350604 351678
rect 386004 351676 386604 351678
rect 422004 351676 422604 351678
rect 458004 351676 458604 351678
rect 494004 351676 494604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 589920 351676 590520 351678
rect -6596 351654 590520 351676
rect -6596 351418 -6414 351654
rect -6178 351418 26186 351654
rect 26422 351418 62186 351654
rect 62422 351418 98186 351654
rect 98422 351418 134186 351654
rect 134422 351418 170186 351654
rect 170422 351418 206186 351654
rect 206422 351418 242186 351654
rect 242422 351418 278186 351654
rect 278422 351418 314186 351654
rect 314422 351418 350186 351654
rect 350422 351418 386186 351654
rect 386422 351418 422186 351654
rect 422422 351418 458186 351654
rect 458422 351418 494186 351654
rect 494422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590102 351654
rect 590338 351418 590520 351654
rect -6596 351334 590520 351418
rect -6596 351098 -6414 351334
rect -6178 351098 26186 351334
rect 26422 351098 62186 351334
rect 62422 351098 98186 351334
rect 98422 351098 134186 351334
rect 134422 351098 170186 351334
rect 170422 351098 206186 351334
rect 206422 351098 242186 351334
rect 242422 351098 278186 351334
rect 278422 351098 314186 351334
rect 314422 351098 350186 351334
rect 350422 351098 386186 351334
rect 386422 351098 422186 351334
rect 422422 351098 458186 351334
rect 458422 351098 494186 351334
rect 494422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590102 351334
rect 590338 351098 590520 351334
rect -6596 351076 590520 351098
rect -6596 351074 -5996 351076
rect 26004 351074 26604 351076
rect 62004 351074 62604 351076
rect 98004 351074 98604 351076
rect 134004 351074 134604 351076
rect 170004 351074 170604 351076
rect 206004 351074 206604 351076
rect 242004 351074 242604 351076
rect 278004 351074 278604 351076
rect 314004 351074 314604 351076
rect 350004 351074 350604 351076
rect 386004 351074 386604 351076
rect 422004 351074 422604 351076
rect 458004 351074 458604 351076
rect 494004 351074 494604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 589920 351074 590520 351076
rect -4756 348076 -4156 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 94404 348076 95004 348078
rect 130404 348076 131004 348078
rect 166404 348076 167004 348078
rect 202404 348076 203004 348078
rect 238404 348076 239004 348078
rect 274404 348076 275004 348078
rect 310404 348076 311004 348078
rect 346404 348076 347004 348078
rect 382404 348076 383004 348078
rect 418404 348076 419004 348078
rect 454404 348076 455004 348078
rect 490404 348076 491004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588080 348076 588680 348078
rect -4756 348054 588680 348076
rect -4756 347818 -4574 348054
rect -4338 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 94586 348054
rect 94822 347818 130586 348054
rect 130822 347818 166586 348054
rect 166822 347818 202586 348054
rect 202822 347818 238586 348054
rect 238822 347818 274586 348054
rect 274822 347818 310586 348054
rect 310822 347818 346586 348054
rect 346822 347818 382586 348054
rect 382822 347818 418586 348054
rect 418822 347818 454586 348054
rect 454822 347818 490586 348054
rect 490822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588262 348054
rect 588498 347818 588680 348054
rect -4756 347734 588680 347818
rect -4756 347498 -4574 347734
rect -4338 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 94586 347734
rect 94822 347498 130586 347734
rect 130822 347498 166586 347734
rect 166822 347498 202586 347734
rect 202822 347498 238586 347734
rect 238822 347498 274586 347734
rect 274822 347498 310586 347734
rect 310822 347498 346586 347734
rect 346822 347498 382586 347734
rect 382822 347498 418586 347734
rect 418822 347498 454586 347734
rect 454822 347498 490586 347734
rect 490822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588262 347734
rect 588498 347498 588680 347734
rect -4756 347476 588680 347498
rect -4756 347474 -4156 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 94404 347474 95004 347476
rect 130404 347474 131004 347476
rect 166404 347474 167004 347476
rect 202404 347474 203004 347476
rect 238404 347474 239004 347476
rect 274404 347474 275004 347476
rect 310404 347474 311004 347476
rect 346404 347474 347004 347476
rect 382404 347474 383004 347476
rect 418404 347474 419004 347476
rect 454404 347474 455004 347476
rect 490404 347474 491004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588080 347474 588680 347476
rect -2916 344476 -2316 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 90804 344476 91404 344478
rect 126804 344476 127404 344478
rect 162804 344476 163404 344478
rect 198804 344476 199404 344478
rect 234804 344476 235404 344478
rect 270804 344476 271404 344478
rect 306804 344476 307404 344478
rect 342804 344476 343404 344478
rect 378804 344476 379404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586240 344476 586840 344478
rect -2916 344454 586840 344476
rect -2916 344218 -2734 344454
rect -2498 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 162986 344454
rect 163222 344218 198986 344454
rect 199222 344218 234986 344454
rect 235222 344218 270986 344454
rect 271222 344218 306986 344454
rect 307222 344218 342986 344454
rect 343222 344218 378986 344454
rect 379222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586422 344454
rect 586658 344218 586840 344454
rect -2916 344134 586840 344218
rect -2916 343898 -2734 344134
rect -2498 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 162986 344134
rect 163222 343898 198986 344134
rect 199222 343898 234986 344134
rect 235222 343898 270986 344134
rect 271222 343898 306986 344134
rect 307222 343898 342986 344134
rect 343222 343898 378986 344134
rect 379222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586422 344134
rect 586658 343898 586840 344134
rect -2916 343876 586840 343898
rect -2916 343874 -2316 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 90804 343874 91404 343876
rect 126804 343874 127404 343876
rect 162804 343874 163404 343876
rect 198804 343874 199404 343876
rect 234804 343874 235404 343876
rect 270804 343874 271404 343876
rect 306804 343874 307404 343876
rect 342804 343874 343404 343876
rect 378804 343874 379404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586240 343874 586840 343876
rect -7516 337276 -6916 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 83604 337276 84204 337278
rect 119604 337276 120204 337278
rect 155604 337276 156204 337278
rect 191604 337276 192204 337278
rect 227604 337276 228204 337278
rect 263604 337276 264204 337278
rect 299604 337276 300204 337278
rect 335604 337276 336204 337278
rect 371604 337276 372204 337278
rect 407604 337276 408204 337278
rect 443604 337276 444204 337278
rect 479604 337276 480204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590840 337276 591440 337278
rect -8436 337254 592360 337276
rect -8436 337018 -7334 337254
rect -7098 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 83786 337254
rect 84022 337018 119786 337254
rect 120022 337018 155786 337254
rect 156022 337018 191786 337254
rect 192022 337018 227786 337254
rect 228022 337018 263786 337254
rect 264022 337018 299786 337254
rect 300022 337018 335786 337254
rect 336022 337018 371786 337254
rect 372022 337018 407786 337254
rect 408022 337018 443786 337254
rect 444022 337018 479786 337254
rect 480022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591022 337254
rect 591258 337018 592360 337254
rect -8436 336934 592360 337018
rect -8436 336698 -7334 336934
rect -7098 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 83786 336934
rect 84022 336698 119786 336934
rect 120022 336698 155786 336934
rect 156022 336698 191786 336934
rect 192022 336698 227786 336934
rect 228022 336698 263786 336934
rect 264022 336698 299786 336934
rect 300022 336698 335786 336934
rect 336022 336698 371786 336934
rect 372022 336698 407786 336934
rect 408022 336698 443786 336934
rect 444022 336698 479786 336934
rect 480022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591022 336934
rect 591258 336698 592360 336934
rect -8436 336676 592360 336698
rect -7516 336674 -6916 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 83604 336674 84204 336676
rect 119604 336674 120204 336676
rect 155604 336674 156204 336676
rect 191604 336674 192204 336676
rect 227604 336674 228204 336676
rect 263604 336674 264204 336676
rect 299604 336674 300204 336676
rect 335604 336674 336204 336676
rect 371604 336674 372204 336676
rect 407604 336674 408204 336676
rect 443604 336674 444204 336676
rect 479604 336674 480204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590840 336674 591440 336676
rect -5676 333676 -5076 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 80004 333676 80604 333678
rect 116004 333676 116604 333678
rect 152004 333676 152604 333678
rect 188004 333676 188604 333678
rect 224004 333676 224604 333678
rect 260004 333676 260604 333678
rect 296004 333676 296604 333678
rect 332004 333676 332604 333678
rect 368004 333676 368604 333678
rect 404004 333676 404604 333678
rect 440004 333676 440604 333678
rect 476004 333676 476604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589000 333676 589600 333678
rect -6596 333654 590520 333676
rect -6596 333418 -5494 333654
rect -5258 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 80186 333654
rect 80422 333418 116186 333654
rect 116422 333418 152186 333654
rect 152422 333418 188186 333654
rect 188422 333418 224186 333654
rect 224422 333418 260186 333654
rect 260422 333418 296186 333654
rect 296422 333418 332186 333654
rect 332422 333418 368186 333654
rect 368422 333418 404186 333654
rect 404422 333418 440186 333654
rect 440422 333418 476186 333654
rect 476422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589182 333654
rect 589418 333418 590520 333654
rect -6596 333334 590520 333418
rect -6596 333098 -5494 333334
rect -5258 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 80186 333334
rect 80422 333098 116186 333334
rect 116422 333098 152186 333334
rect 152422 333098 188186 333334
rect 188422 333098 224186 333334
rect 224422 333098 260186 333334
rect 260422 333098 296186 333334
rect 296422 333098 332186 333334
rect 332422 333098 368186 333334
rect 368422 333098 404186 333334
rect 404422 333098 440186 333334
rect 440422 333098 476186 333334
rect 476422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589182 333334
rect 589418 333098 590520 333334
rect -6596 333076 590520 333098
rect -5676 333074 -5076 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 80004 333074 80604 333076
rect 116004 333074 116604 333076
rect 152004 333074 152604 333076
rect 188004 333074 188604 333076
rect 224004 333074 224604 333076
rect 260004 333074 260604 333076
rect 296004 333074 296604 333076
rect 332004 333074 332604 333076
rect 368004 333074 368604 333076
rect 404004 333074 404604 333076
rect 440004 333074 440604 333076
rect 476004 333074 476604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589000 333074 589600 333076
rect -3836 330076 -3236 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 112404 330076 113004 330078
rect 148404 330076 149004 330078
rect 184404 330076 185004 330078
rect 220404 330076 221004 330078
rect 256404 330076 257004 330078
rect 292404 330076 293004 330078
rect 328404 330076 329004 330078
rect 364404 330076 365004 330078
rect 400404 330076 401004 330078
rect 436404 330076 437004 330078
rect 472404 330076 473004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587160 330076 587760 330078
rect -4756 330054 588680 330076
rect -4756 329818 -3654 330054
rect -3418 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 112586 330054
rect 112822 329818 148586 330054
rect 148822 329818 184586 330054
rect 184822 329818 220586 330054
rect 220822 329818 256586 330054
rect 256822 329818 292586 330054
rect 292822 329818 328586 330054
rect 328822 329818 364586 330054
rect 364822 329818 400586 330054
rect 400822 329818 436586 330054
rect 436822 329818 472586 330054
rect 472822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587342 330054
rect 587578 329818 588680 330054
rect -4756 329734 588680 329818
rect -4756 329498 -3654 329734
rect -3418 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 112586 329734
rect 112822 329498 148586 329734
rect 148822 329498 184586 329734
rect 184822 329498 220586 329734
rect 220822 329498 256586 329734
rect 256822 329498 292586 329734
rect 292822 329498 328586 329734
rect 328822 329498 364586 329734
rect 364822 329498 400586 329734
rect 400822 329498 436586 329734
rect 436822 329498 472586 329734
rect 472822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587342 329734
rect 587578 329498 588680 329734
rect -4756 329476 588680 329498
rect -3836 329474 -3236 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 112404 329474 113004 329476
rect 148404 329474 149004 329476
rect 184404 329474 185004 329476
rect 220404 329474 221004 329476
rect 256404 329474 257004 329476
rect 292404 329474 293004 329476
rect 328404 329474 329004 329476
rect 364404 329474 365004 329476
rect 400404 329474 401004 329476
rect 436404 329474 437004 329476
rect 472404 329474 473004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587160 329474 587760 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 144804 326476 145404 326478
rect 180804 326476 181404 326478
rect 216804 326476 217404 326478
rect 252804 326476 253404 326478
rect 288804 326476 289404 326478
rect 324804 326476 325404 326478
rect 360804 326476 361404 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2916 326454 586840 326476
rect -2916 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 180986 326454
rect 181222 326218 216986 326454
rect 217222 326218 252986 326454
rect 253222 326218 288986 326454
rect 289222 326218 324986 326454
rect 325222 326218 360986 326454
rect 361222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586840 326454
rect -2916 326134 586840 326218
rect -2916 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 180986 326134
rect 181222 325898 216986 326134
rect 217222 325898 252986 326134
rect 253222 325898 288986 326134
rect 289222 325898 324986 326134
rect 325222 325898 360986 326134
rect 361222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586840 326134
rect -2916 325876 586840 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 144804 325874 145404 325876
rect 180804 325874 181404 325876
rect 216804 325874 217404 325876
rect 252804 325874 253404 325876
rect 288804 325874 289404 325876
rect 324804 325874 325404 325876
rect 360804 325874 361404 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8436 319276 -7836 319278
rect 29604 319276 30204 319278
rect 65604 319276 66204 319278
rect 101604 319276 102204 319278
rect 137604 319276 138204 319278
rect 173604 319276 174204 319278
rect 209604 319276 210204 319278
rect 245604 319276 246204 319278
rect 281604 319276 282204 319278
rect 317604 319276 318204 319278
rect 353604 319276 354204 319278
rect 389604 319276 390204 319278
rect 425604 319276 426204 319278
rect 461604 319276 462204 319278
rect 497604 319276 498204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591760 319276 592360 319278
rect -8436 319254 592360 319276
rect -8436 319018 -8254 319254
rect -8018 319018 29786 319254
rect 30022 319018 65786 319254
rect 66022 319018 101786 319254
rect 102022 319018 137786 319254
rect 138022 319018 173786 319254
rect 174022 319018 209786 319254
rect 210022 319018 245786 319254
rect 246022 319018 281786 319254
rect 282022 319018 317786 319254
rect 318022 319018 353786 319254
rect 354022 319018 389786 319254
rect 390022 319018 425786 319254
rect 426022 319018 461786 319254
rect 462022 319018 497786 319254
rect 498022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 591942 319254
rect 592178 319018 592360 319254
rect -8436 318934 592360 319018
rect -8436 318698 -8254 318934
rect -8018 318698 29786 318934
rect 30022 318698 65786 318934
rect 66022 318698 101786 318934
rect 102022 318698 137786 318934
rect 138022 318698 173786 318934
rect 174022 318698 209786 318934
rect 210022 318698 245786 318934
rect 246022 318698 281786 318934
rect 282022 318698 317786 318934
rect 318022 318698 353786 318934
rect 354022 318698 389786 318934
rect 390022 318698 425786 318934
rect 426022 318698 461786 318934
rect 462022 318698 497786 318934
rect 498022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 591942 318934
rect 592178 318698 592360 318934
rect -8436 318676 592360 318698
rect -8436 318674 -7836 318676
rect 29604 318674 30204 318676
rect 65604 318674 66204 318676
rect 101604 318674 102204 318676
rect 137604 318674 138204 318676
rect 173604 318674 174204 318676
rect 209604 318674 210204 318676
rect 245604 318674 246204 318676
rect 281604 318674 282204 318676
rect 317604 318674 318204 318676
rect 353604 318674 354204 318676
rect 389604 318674 390204 318676
rect 425604 318674 426204 318676
rect 461604 318674 462204 318676
rect 497604 318674 498204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591760 318674 592360 318676
rect -6596 315676 -5996 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 98004 315676 98604 315678
rect 134004 315676 134604 315678
rect 170004 315676 170604 315678
rect 206004 315676 206604 315678
rect 242004 315676 242604 315678
rect 278004 315676 278604 315678
rect 314004 315676 314604 315678
rect 350004 315676 350604 315678
rect 386004 315676 386604 315678
rect 422004 315676 422604 315678
rect 458004 315676 458604 315678
rect 494004 315676 494604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 589920 315676 590520 315678
rect -6596 315654 590520 315676
rect -6596 315418 -6414 315654
rect -6178 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 98186 315654
rect 98422 315418 134186 315654
rect 134422 315418 170186 315654
rect 170422 315418 206186 315654
rect 206422 315418 242186 315654
rect 242422 315418 278186 315654
rect 278422 315418 314186 315654
rect 314422 315418 350186 315654
rect 350422 315418 386186 315654
rect 386422 315418 422186 315654
rect 422422 315418 458186 315654
rect 458422 315418 494186 315654
rect 494422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590102 315654
rect 590338 315418 590520 315654
rect -6596 315334 590520 315418
rect -6596 315098 -6414 315334
rect -6178 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 98186 315334
rect 98422 315098 134186 315334
rect 134422 315098 170186 315334
rect 170422 315098 206186 315334
rect 206422 315098 242186 315334
rect 242422 315098 278186 315334
rect 278422 315098 314186 315334
rect 314422 315098 350186 315334
rect 350422 315098 386186 315334
rect 386422 315098 422186 315334
rect 422422 315098 458186 315334
rect 458422 315098 494186 315334
rect 494422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590102 315334
rect 590338 315098 590520 315334
rect -6596 315076 590520 315098
rect -6596 315074 -5996 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 98004 315074 98604 315076
rect 134004 315074 134604 315076
rect 170004 315074 170604 315076
rect 206004 315074 206604 315076
rect 242004 315074 242604 315076
rect 278004 315074 278604 315076
rect 314004 315074 314604 315076
rect 350004 315074 350604 315076
rect 386004 315074 386604 315076
rect 422004 315074 422604 315076
rect 458004 315074 458604 315076
rect 494004 315074 494604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 589920 315074 590520 315076
rect -4756 312076 -4156 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 94404 312076 95004 312078
rect 130404 312076 131004 312078
rect 166404 312076 167004 312078
rect 202404 312076 203004 312078
rect 238404 312076 239004 312078
rect 274404 312076 275004 312078
rect 310404 312076 311004 312078
rect 346404 312076 347004 312078
rect 382404 312076 383004 312078
rect 418404 312076 419004 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588080 312076 588680 312078
rect -4756 312054 588680 312076
rect -4756 311818 -4574 312054
rect -4338 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 94586 312054
rect 94822 311818 130586 312054
rect 130822 311818 166586 312054
rect 166822 311818 202586 312054
rect 202822 311818 238586 312054
rect 238822 311818 274586 312054
rect 274822 311818 310586 312054
rect 310822 311818 346586 312054
rect 346822 311818 382586 312054
rect 382822 311818 418586 312054
rect 418822 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588262 312054
rect 588498 311818 588680 312054
rect -4756 311734 588680 311818
rect -4756 311498 -4574 311734
rect -4338 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 94586 311734
rect 94822 311498 130586 311734
rect 130822 311498 166586 311734
rect 166822 311498 202586 311734
rect 202822 311498 238586 311734
rect 238822 311498 274586 311734
rect 274822 311498 310586 311734
rect 310822 311498 346586 311734
rect 346822 311498 382586 311734
rect 382822 311498 418586 311734
rect 418822 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588262 311734
rect 588498 311498 588680 311734
rect -4756 311476 588680 311498
rect -4756 311474 -4156 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 94404 311474 95004 311476
rect 130404 311474 131004 311476
rect 166404 311474 167004 311476
rect 202404 311474 203004 311476
rect 238404 311474 239004 311476
rect 274404 311474 275004 311476
rect 310404 311474 311004 311476
rect 346404 311474 347004 311476
rect 382404 311474 383004 311476
rect 418404 311474 419004 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588080 311474 588680 311476
rect -2916 308476 -2316 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 270804 308476 271404 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586240 308476 586840 308478
rect -2916 308454 586840 308476
rect -2916 308218 -2734 308454
rect -2498 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586422 308454
rect 586658 308218 586840 308454
rect -2916 308134 586840 308218
rect -2916 307898 -2734 308134
rect -2498 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586422 308134
rect 586658 307898 586840 308134
rect -2916 307876 586840 307898
rect -2916 307874 -2316 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 270804 307874 271404 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586240 307874 586840 307876
rect -7516 301276 -6916 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 83604 301276 84204 301278
rect 119604 301276 120204 301278
rect 155604 301276 156204 301278
rect 191604 301276 192204 301278
rect 227604 301276 228204 301278
rect 263604 301276 264204 301278
rect 299604 301276 300204 301278
rect 335604 301276 336204 301278
rect 371604 301276 372204 301278
rect 407604 301276 408204 301278
rect 443604 301276 444204 301278
rect 479604 301276 480204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590840 301276 591440 301278
rect -8436 301254 592360 301276
rect -8436 301018 -7334 301254
rect -7098 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 83786 301254
rect 84022 301018 119786 301254
rect 120022 301018 155786 301254
rect 156022 301018 191786 301254
rect 192022 301018 227786 301254
rect 228022 301018 263786 301254
rect 264022 301018 299786 301254
rect 300022 301018 335786 301254
rect 336022 301018 371786 301254
rect 372022 301018 407786 301254
rect 408022 301018 443786 301254
rect 444022 301018 479786 301254
rect 480022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591022 301254
rect 591258 301018 592360 301254
rect -8436 300934 592360 301018
rect -8436 300698 -7334 300934
rect -7098 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 83786 300934
rect 84022 300698 119786 300934
rect 120022 300698 155786 300934
rect 156022 300698 191786 300934
rect 192022 300698 227786 300934
rect 228022 300698 263786 300934
rect 264022 300698 299786 300934
rect 300022 300698 335786 300934
rect 336022 300698 371786 300934
rect 372022 300698 407786 300934
rect 408022 300698 443786 300934
rect 444022 300698 479786 300934
rect 480022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591022 300934
rect 591258 300698 592360 300934
rect -8436 300676 592360 300698
rect -7516 300674 -6916 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 83604 300674 84204 300676
rect 119604 300674 120204 300676
rect 155604 300674 156204 300676
rect 191604 300674 192204 300676
rect 227604 300674 228204 300676
rect 263604 300674 264204 300676
rect 299604 300674 300204 300676
rect 335604 300674 336204 300676
rect 371604 300674 372204 300676
rect 407604 300674 408204 300676
rect 443604 300674 444204 300676
rect 479604 300674 480204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590840 300674 591440 300676
rect -5676 297676 -5076 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 116004 297676 116604 297678
rect 152004 297676 152604 297678
rect 188004 297676 188604 297678
rect 224004 297676 224604 297678
rect 260004 297676 260604 297678
rect 296004 297676 296604 297678
rect 332004 297676 332604 297678
rect 368004 297676 368604 297678
rect 404004 297676 404604 297678
rect 440004 297676 440604 297678
rect 476004 297676 476604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589000 297676 589600 297678
rect -6596 297654 590520 297676
rect -6596 297418 -5494 297654
rect -5258 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 116186 297654
rect 116422 297418 152186 297654
rect 152422 297418 188186 297654
rect 188422 297418 224186 297654
rect 224422 297418 260186 297654
rect 260422 297418 296186 297654
rect 296422 297418 332186 297654
rect 332422 297418 368186 297654
rect 368422 297418 404186 297654
rect 404422 297418 440186 297654
rect 440422 297418 476186 297654
rect 476422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589182 297654
rect 589418 297418 590520 297654
rect -6596 297334 590520 297418
rect -6596 297098 -5494 297334
rect -5258 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 116186 297334
rect 116422 297098 152186 297334
rect 152422 297098 188186 297334
rect 188422 297098 224186 297334
rect 224422 297098 260186 297334
rect 260422 297098 296186 297334
rect 296422 297098 332186 297334
rect 332422 297098 368186 297334
rect 368422 297098 404186 297334
rect 404422 297098 440186 297334
rect 440422 297098 476186 297334
rect 476422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589182 297334
rect 589418 297098 590520 297334
rect -6596 297076 590520 297098
rect -5676 297074 -5076 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 116004 297074 116604 297076
rect 152004 297074 152604 297076
rect 188004 297074 188604 297076
rect 224004 297074 224604 297076
rect 260004 297074 260604 297076
rect 296004 297074 296604 297076
rect 332004 297074 332604 297076
rect 368004 297074 368604 297076
rect 404004 297074 404604 297076
rect 440004 297074 440604 297076
rect 476004 297074 476604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589000 297074 589600 297076
rect -3836 294076 -3236 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 148404 294076 149004 294078
rect 184404 294076 185004 294078
rect 220404 294076 221004 294078
rect 256404 294076 257004 294078
rect 292404 294076 293004 294078
rect 328404 294076 329004 294078
rect 364404 294076 365004 294078
rect 400404 294076 401004 294078
rect 436404 294076 437004 294078
rect 472404 294076 473004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587160 294076 587760 294078
rect -4756 294054 588680 294076
rect -4756 293818 -3654 294054
rect -3418 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 148586 294054
rect 148822 293818 184586 294054
rect 184822 293818 220586 294054
rect 220822 293818 256586 294054
rect 256822 293818 292586 294054
rect 292822 293818 328586 294054
rect 328822 293818 364586 294054
rect 364822 293818 400586 294054
rect 400822 293818 436586 294054
rect 436822 293818 472586 294054
rect 472822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587342 294054
rect 587578 293818 588680 294054
rect -4756 293734 588680 293818
rect -4756 293498 -3654 293734
rect -3418 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 148586 293734
rect 148822 293498 184586 293734
rect 184822 293498 220586 293734
rect 220822 293498 256586 293734
rect 256822 293498 292586 293734
rect 292822 293498 328586 293734
rect 328822 293498 364586 293734
rect 364822 293498 400586 293734
rect 400822 293498 436586 293734
rect 436822 293498 472586 293734
rect 472822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587342 293734
rect 587578 293498 588680 293734
rect -4756 293476 588680 293498
rect -3836 293474 -3236 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 148404 293474 149004 293476
rect 184404 293474 185004 293476
rect 220404 293474 221004 293476
rect 256404 293474 257004 293476
rect 292404 293474 293004 293476
rect 328404 293474 329004 293476
rect 364404 293474 365004 293476
rect 400404 293474 401004 293476
rect 436404 293474 437004 293476
rect 472404 293474 473004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587160 293474 587760 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 288804 290476 289404 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2916 290454 586840 290476
rect -2916 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586840 290454
rect -2916 290134 586840 290218
rect -2916 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586840 290134
rect -2916 289876 586840 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 288804 289874 289404 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8436 283276 -7836 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 101604 283276 102204 283278
rect 137604 283276 138204 283278
rect 173604 283276 174204 283278
rect 209604 283276 210204 283278
rect 245604 283276 246204 283278
rect 281604 283276 282204 283278
rect 317604 283276 318204 283278
rect 353604 283276 354204 283278
rect 389604 283276 390204 283278
rect 425604 283276 426204 283278
rect 461604 283276 462204 283278
rect 497604 283276 498204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591760 283276 592360 283278
rect -8436 283254 592360 283276
rect -8436 283018 -8254 283254
rect -8018 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 101786 283254
rect 102022 283018 137786 283254
rect 138022 283018 173786 283254
rect 174022 283018 209786 283254
rect 210022 283018 245786 283254
rect 246022 283018 281786 283254
rect 282022 283018 317786 283254
rect 318022 283018 353786 283254
rect 354022 283018 389786 283254
rect 390022 283018 425786 283254
rect 426022 283018 461786 283254
rect 462022 283018 497786 283254
rect 498022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 591942 283254
rect 592178 283018 592360 283254
rect -8436 282934 592360 283018
rect -8436 282698 -8254 282934
rect -8018 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 101786 282934
rect 102022 282698 137786 282934
rect 138022 282698 173786 282934
rect 174022 282698 209786 282934
rect 210022 282698 245786 282934
rect 246022 282698 281786 282934
rect 282022 282698 317786 282934
rect 318022 282698 353786 282934
rect 354022 282698 389786 282934
rect 390022 282698 425786 282934
rect 426022 282698 461786 282934
rect 462022 282698 497786 282934
rect 498022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 591942 282934
rect 592178 282698 592360 282934
rect -8436 282676 592360 282698
rect -8436 282674 -7836 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 101604 282674 102204 282676
rect 137604 282674 138204 282676
rect 173604 282674 174204 282676
rect 209604 282674 210204 282676
rect 245604 282674 246204 282676
rect 281604 282674 282204 282676
rect 317604 282674 318204 282676
rect 353604 282674 354204 282676
rect 389604 282674 390204 282676
rect 425604 282674 426204 282676
rect 461604 282674 462204 282676
rect 497604 282674 498204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591760 282674 592360 282676
rect -6596 279676 -5996 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 98004 279676 98604 279678
rect 134004 279676 134604 279678
rect 170004 279676 170604 279678
rect 206004 279676 206604 279678
rect 242004 279676 242604 279678
rect 278004 279676 278604 279678
rect 314004 279676 314604 279678
rect 350004 279676 350604 279678
rect 386004 279676 386604 279678
rect 422004 279676 422604 279678
rect 458004 279676 458604 279678
rect 494004 279676 494604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 589920 279676 590520 279678
rect -6596 279654 590520 279676
rect -6596 279418 -6414 279654
rect -6178 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 98186 279654
rect 98422 279418 134186 279654
rect 134422 279418 170186 279654
rect 170422 279418 206186 279654
rect 206422 279418 242186 279654
rect 242422 279418 278186 279654
rect 278422 279418 314186 279654
rect 314422 279418 350186 279654
rect 350422 279418 386186 279654
rect 386422 279418 422186 279654
rect 422422 279418 458186 279654
rect 458422 279418 494186 279654
rect 494422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590102 279654
rect 590338 279418 590520 279654
rect -6596 279334 590520 279418
rect -6596 279098 -6414 279334
rect -6178 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 98186 279334
rect 98422 279098 134186 279334
rect 134422 279098 170186 279334
rect 170422 279098 206186 279334
rect 206422 279098 242186 279334
rect 242422 279098 278186 279334
rect 278422 279098 314186 279334
rect 314422 279098 350186 279334
rect 350422 279098 386186 279334
rect 386422 279098 422186 279334
rect 422422 279098 458186 279334
rect 458422 279098 494186 279334
rect 494422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590102 279334
rect 590338 279098 590520 279334
rect -6596 279076 590520 279098
rect -6596 279074 -5996 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 98004 279074 98604 279076
rect 134004 279074 134604 279076
rect 170004 279074 170604 279076
rect 206004 279074 206604 279076
rect 242004 279074 242604 279076
rect 278004 279074 278604 279076
rect 314004 279074 314604 279076
rect 350004 279074 350604 279076
rect 386004 279074 386604 279076
rect 422004 279074 422604 279076
rect 458004 279074 458604 279076
rect 494004 279074 494604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 589920 279074 590520 279076
rect -4756 276076 -4156 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 166404 276076 167004 276078
rect 202404 276076 203004 276078
rect 238404 276076 239004 276078
rect 274404 276076 275004 276078
rect 310404 276076 311004 276078
rect 346404 276076 347004 276078
rect 382404 276076 383004 276078
rect 418404 276076 419004 276078
rect 454404 276076 455004 276078
rect 490404 276076 491004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588080 276076 588680 276078
rect -4756 276054 588680 276076
rect -4756 275818 -4574 276054
rect -4338 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 166586 276054
rect 166822 275818 202586 276054
rect 202822 275818 238586 276054
rect 238822 275818 274586 276054
rect 274822 275818 310586 276054
rect 310822 275818 346586 276054
rect 346822 275818 382586 276054
rect 382822 275818 418586 276054
rect 418822 275818 454586 276054
rect 454822 275818 490586 276054
rect 490822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588262 276054
rect 588498 275818 588680 276054
rect -4756 275734 588680 275818
rect -4756 275498 -4574 275734
rect -4338 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 166586 275734
rect 166822 275498 202586 275734
rect 202822 275498 238586 275734
rect 238822 275498 274586 275734
rect 274822 275498 310586 275734
rect 310822 275498 346586 275734
rect 346822 275498 382586 275734
rect 382822 275498 418586 275734
rect 418822 275498 454586 275734
rect 454822 275498 490586 275734
rect 490822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588262 275734
rect 588498 275498 588680 275734
rect -4756 275476 588680 275498
rect -4756 275474 -4156 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 166404 275474 167004 275476
rect 202404 275474 203004 275476
rect 238404 275474 239004 275476
rect 274404 275474 275004 275476
rect 310404 275474 311004 275476
rect 346404 275474 347004 275476
rect 382404 275474 383004 275476
rect 418404 275474 419004 275476
rect 454404 275474 455004 275476
rect 490404 275474 491004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588080 275474 588680 275476
rect -2916 272476 -2316 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 198804 272476 199404 272478
rect 234804 272476 235404 272478
rect 270804 272476 271404 272478
rect 306804 272476 307404 272478
rect 342804 272476 343404 272478
rect 378804 272476 379404 272478
rect 414804 272476 415404 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586240 272476 586840 272478
rect -2916 272454 586840 272476
rect -2916 272218 -2734 272454
rect -2498 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 198986 272454
rect 199222 272218 234986 272454
rect 235222 272218 270986 272454
rect 271222 272218 306986 272454
rect 307222 272218 342986 272454
rect 343222 272218 378986 272454
rect 379222 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586422 272454
rect 586658 272218 586840 272454
rect -2916 272134 586840 272218
rect -2916 271898 -2734 272134
rect -2498 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 198986 272134
rect 199222 271898 234986 272134
rect 235222 271898 270986 272134
rect 271222 271898 306986 272134
rect 307222 271898 342986 272134
rect 343222 271898 378986 272134
rect 379222 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586422 272134
rect 586658 271898 586840 272134
rect -2916 271876 586840 271898
rect -2916 271874 -2316 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 198804 271874 199404 271876
rect 234804 271874 235404 271876
rect 270804 271874 271404 271876
rect 306804 271874 307404 271876
rect 342804 271874 343404 271876
rect 378804 271874 379404 271876
rect 414804 271874 415404 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586240 271874 586840 271876
rect -7516 265276 -6916 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 83604 265276 84204 265278
rect 119604 265276 120204 265278
rect 155604 265276 156204 265278
rect 191604 265276 192204 265278
rect 227604 265276 228204 265278
rect 263604 265276 264204 265278
rect 299604 265276 300204 265278
rect 335604 265276 336204 265278
rect 371604 265276 372204 265278
rect 407604 265276 408204 265278
rect 443604 265276 444204 265278
rect 479604 265276 480204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590840 265276 591440 265278
rect -8436 265254 592360 265276
rect -8436 265018 -7334 265254
rect -7098 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 83786 265254
rect 84022 265018 119786 265254
rect 120022 265018 155786 265254
rect 156022 265018 191786 265254
rect 192022 265018 227786 265254
rect 228022 265018 263786 265254
rect 264022 265018 299786 265254
rect 300022 265018 335786 265254
rect 336022 265018 371786 265254
rect 372022 265018 407786 265254
rect 408022 265018 443786 265254
rect 444022 265018 479786 265254
rect 480022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591022 265254
rect 591258 265018 592360 265254
rect -8436 264934 592360 265018
rect -8436 264698 -7334 264934
rect -7098 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 83786 264934
rect 84022 264698 119786 264934
rect 120022 264698 155786 264934
rect 156022 264698 191786 264934
rect 192022 264698 227786 264934
rect 228022 264698 263786 264934
rect 264022 264698 299786 264934
rect 300022 264698 335786 264934
rect 336022 264698 371786 264934
rect 372022 264698 407786 264934
rect 408022 264698 443786 264934
rect 444022 264698 479786 264934
rect 480022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591022 264934
rect 591258 264698 592360 264934
rect -8436 264676 592360 264698
rect -7516 264674 -6916 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 83604 264674 84204 264676
rect 119604 264674 120204 264676
rect 155604 264674 156204 264676
rect 191604 264674 192204 264676
rect 227604 264674 228204 264676
rect 263604 264674 264204 264676
rect 299604 264674 300204 264676
rect 335604 264674 336204 264676
rect 371604 264674 372204 264676
rect 407604 264674 408204 264676
rect 443604 264674 444204 264676
rect 479604 264674 480204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590840 264674 591440 264676
rect -5676 261676 -5076 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 116004 261676 116604 261678
rect 152004 261676 152604 261678
rect 188004 261676 188604 261678
rect 224004 261676 224604 261678
rect 260004 261676 260604 261678
rect 296004 261676 296604 261678
rect 332004 261676 332604 261678
rect 368004 261676 368604 261678
rect 404004 261676 404604 261678
rect 440004 261676 440604 261678
rect 476004 261676 476604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589000 261676 589600 261678
rect -6596 261654 590520 261676
rect -6596 261418 -5494 261654
rect -5258 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 116186 261654
rect 116422 261418 152186 261654
rect 152422 261418 188186 261654
rect 188422 261418 224186 261654
rect 224422 261418 260186 261654
rect 260422 261418 296186 261654
rect 296422 261418 332186 261654
rect 332422 261418 368186 261654
rect 368422 261418 404186 261654
rect 404422 261418 440186 261654
rect 440422 261418 476186 261654
rect 476422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589182 261654
rect 589418 261418 590520 261654
rect -6596 261334 590520 261418
rect -6596 261098 -5494 261334
rect -5258 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 116186 261334
rect 116422 261098 152186 261334
rect 152422 261098 188186 261334
rect 188422 261098 224186 261334
rect 224422 261098 260186 261334
rect 260422 261098 296186 261334
rect 296422 261098 332186 261334
rect 332422 261098 368186 261334
rect 368422 261098 404186 261334
rect 404422 261098 440186 261334
rect 440422 261098 476186 261334
rect 476422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589182 261334
rect 589418 261098 590520 261334
rect -6596 261076 590520 261098
rect -5676 261074 -5076 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 116004 261074 116604 261076
rect 152004 261074 152604 261076
rect 188004 261074 188604 261076
rect 224004 261074 224604 261076
rect 260004 261074 260604 261076
rect 296004 261074 296604 261076
rect 332004 261074 332604 261076
rect 368004 261074 368604 261076
rect 404004 261074 404604 261076
rect 440004 261074 440604 261076
rect 476004 261074 476604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589000 261074 589600 261076
rect -3836 258076 -3236 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 148404 258076 149004 258078
rect 184404 258076 185004 258078
rect 220404 258076 221004 258078
rect 256404 258076 257004 258078
rect 292404 258076 293004 258078
rect 328404 258076 329004 258078
rect 364404 258076 365004 258078
rect 400404 258076 401004 258078
rect 436404 258076 437004 258078
rect 472404 258076 473004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587160 258076 587760 258078
rect -4756 258054 588680 258076
rect -4756 257818 -3654 258054
rect -3418 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 148586 258054
rect 148822 257818 184586 258054
rect 184822 257818 220586 258054
rect 220822 257818 256586 258054
rect 256822 257818 292586 258054
rect 292822 257818 328586 258054
rect 328822 257818 364586 258054
rect 364822 257818 400586 258054
rect 400822 257818 436586 258054
rect 436822 257818 472586 258054
rect 472822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587342 258054
rect 587578 257818 588680 258054
rect -4756 257734 588680 257818
rect -4756 257498 -3654 257734
rect -3418 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 148586 257734
rect 148822 257498 184586 257734
rect 184822 257498 220586 257734
rect 220822 257498 256586 257734
rect 256822 257498 292586 257734
rect 292822 257498 328586 257734
rect 328822 257498 364586 257734
rect 364822 257498 400586 257734
rect 400822 257498 436586 257734
rect 436822 257498 472586 257734
rect 472822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587342 257734
rect 587578 257498 588680 257734
rect -4756 257476 588680 257498
rect -3836 257474 -3236 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 148404 257474 149004 257476
rect 184404 257474 185004 257476
rect 220404 257474 221004 257476
rect 256404 257474 257004 257476
rect 292404 257474 293004 257476
rect 328404 257474 329004 257476
rect 364404 257474 365004 257476
rect 400404 257474 401004 257476
rect 436404 257474 437004 257476
rect 472404 257474 473004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587160 257474 587760 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 144804 254476 145404 254478
rect 180804 254476 181404 254478
rect 216804 254476 217404 254478
rect 252804 254476 253404 254478
rect 288804 254476 289404 254478
rect 324804 254476 325404 254478
rect 360804 254476 361404 254478
rect 396804 254476 397404 254478
rect 432804 254476 433404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2916 254454 586840 254476
rect -2916 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 216986 254454
rect 217222 254218 252986 254454
rect 253222 254218 288986 254454
rect 289222 254218 324986 254454
rect 325222 254218 360986 254454
rect 361222 254218 396986 254454
rect 397222 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586840 254454
rect -2916 254134 586840 254218
rect -2916 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 216986 254134
rect 217222 253898 252986 254134
rect 253222 253898 288986 254134
rect 289222 253898 324986 254134
rect 325222 253898 360986 254134
rect 361222 253898 396986 254134
rect 397222 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586840 254134
rect -2916 253876 586840 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 144804 253874 145404 253876
rect 180804 253874 181404 253876
rect 216804 253874 217404 253876
rect 252804 253874 253404 253876
rect 288804 253874 289404 253876
rect 324804 253874 325404 253876
rect 360804 253874 361404 253876
rect 396804 253874 397404 253876
rect 432804 253874 433404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8436 247276 -7836 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 101604 247276 102204 247278
rect 137604 247276 138204 247278
rect 173604 247276 174204 247278
rect 209604 247276 210204 247278
rect 245604 247276 246204 247278
rect 281604 247276 282204 247278
rect 317604 247276 318204 247278
rect 353604 247276 354204 247278
rect 389604 247276 390204 247278
rect 425604 247276 426204 247278
rect 461604 247276 462204 247278
rect 497604 247276 498204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591760 247276 592360 247278
rect -8436 247254 592360 247276
rect -8436 247018 -8254 247254
rect -8018 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 101786 247254
rect 102022 247018 137786 247254
rect 138022 247018 173786 247254
rect 174022 247018 209786 247254
rect 210022 247018 245786 247254
rect 246022 247018 281786 247254
rect 282022 247018 317786 247254
rect 318022 247018 353786 247254
rect 354022 247018 389786 247254
rect 390022 247018 425786 247254
rect 426022 247018 461786 247254
rect 462022 247018 497786 247254
rect 498022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 591942 247254
rect 592178 247018 592360 247254
rect -8436 246934 592360 247018
rect -8436 246698 -8254 246934
rect -8018 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 101786 246934
rect 102022 246698 137786 246934
rect 138022 246698 173786 246934
rect 174022 246698 209786 246934
rect 210022 246698 245786 246934
rect 246022 246698 281786 246934
rect 282022 246698 317786 246934
rect 318022 246698 353786 246934
rect 354022 246698 389786 246934
rect 390022 246698 425786 246934
rect 426022 246698 461786 246934
rect 462022 246698 497786 246934
rect 498022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 591942 246934
rect 592178 246698 592360 246934
rect -8436 246676 592360 246698
rect -8436 246674 -7836 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 101604 246674 102204 246676
rect 137604 246674 138204 246676
rect 173604 246674 174204 246676
rect 209604 246674 210204 246676
rect 245604 246674 246204 246676
rect 281604 246674 282204 246676
rect 317604 246674 318204 246676
rect 353604 246674 354204 246676
rect 389604 246674 390204 246676
rect 425604 246674 426204 246676
rect 461604 246674 462204 246676
rect 497604 246674 498204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591760 246674 592360 246676
rect -6596 243676 -5996 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 98004 243676 98604 243678
rect 134004 243676 134604 243678
rect 170004 243676 170604 243678
rect 206004 243676 206604 243678
rect 242004 243676 242604 243678
rect 278004 243676 278604 243678
rect 314004 243676 314604 243678
rect 350004 243676 350604 243678
rect 386004 243676 386604 243678
rect 422004 243676 422604 243678
rect 458004 243676 458604 243678
rect 494004 243676 494604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 589920 243676 590520 243678
rect -6596 243654 590520 243676
rect -6596 243418 -6414 243654
rect -6178 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 98186 243654
rect 98422 243418 134186 243654
rect 134422 243418 170186 243654
rect 170422 243418 206186 243654
rect 206422 243418 242186 243654
rect 242422 243418 278186 243654
rect 278422 243418 314186 243654
rect 314422 243418 350186 243654
rect 350422 243418 386186 243654
rect 386422 243418 422186 243654
rect 422422 243418 458186 243654
rect 458422 243418 494186 243654
rect 494422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590102 243654
rect 590338 243418 590520 243654
rect -6596 243334 590520 243418
rect -6596 243098 -6414 243334
rect -6178 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 98186 243334
rect 98422 243098 134186 243334
rect 134422 243098 170186 243334
rect 170422 243098 206186 243334
rect 206422 243098 242186 243334
rect 242422 243098 278186 243334
rect 278422 243098 314186 243334
rect 314422 243098 350186 243334
rect 350422 243098 386186 243334
rect 386422 243098 422186 243334
rect 422422 243098 458186 243334
rect 458422 243098 494186 243334
rect 494422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590102 243334
rect 590338 243098 590520 243334
rect -6596 243076 590520 243098
rect -6596 243074 -5996 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 98004 243074 98604 243076
rect 134004 243074 134604 243076
rect 170004 243074 170604 243076
rect 206004 243074 206604 243076
rect 242004 243074 242604 243076
rect 278004 243074 278604 243076
rect 314004 243074 314604 243076
rect 350004 243074 350604 243076
rect 386004 243074 386604 243076
rect 422004 243074 422604 243076
rect 458004 243074 458604 243076
rect 494004 243074 494604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 589920 243074 590520 243076
rect -4756 240076 -4156 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 166404 240076 167004 240078
rect 202404 240076 203004 240078
rect 238404 240076 239004 240078
rect 274404 240076 275004 240078
rect 310404 240076 311004 240078
rect 346404 240076 347004 240078
rect 382404 240076 383004 240078
rect 418404 240076 419004 240078
rect 454404 240076 455004 240078
rect 490404 240076 491004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588080 240076 588680 240078
rect -4756 240054 588680 240076
rect -4756 239818 -4574 240054
rect -4338 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 166586 240054
rect 166822 239818 202586 240054
rect 202822 239818 238586 240054
rect 238822 239818 274586 240054
rect 274822 239818 310586 240054
rect 310822 239818 346586 240054
rect 346822 239818 382586 240054
rect 382822 239818 418586 240054
rect 418822 239818 454586 240054
rect 454822 239818 490586 240054
rect 490822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588262 240054
rect 588498 239818 588680 240054
rect -4756 239734 588680 239818
rect -4756 239498 -4574 239734
rect -4338 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 166586 239734
rect 166822 239498 202586 239734
rect 202822 239498 238586 239734
rect 238822 239498 274586 239734
rect 274822 239498 310586 239734
rect 310822 239498 346586 239734
rect 346822 239498 382586 239734
rect 382822 239498 418586 239734
rect 418822 239498 454586 239734
rect 454822 239498 490586 239734
rect 490822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588262 239734
rect 588498 239498 588680 239734
rect -4756 239476 588680 239498
rect -4756 239474 -4156 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 166404 239474 167004 239476
rect 202404 239474 203004 239476
rect 238404 239474 239004 239476
rect 274404 239474 275004 239476
rect 310404 239474 311004 239476
rect 346404 239474 347004 239476
rect 382404 239474 383004 239476
rect 418404 239474 419004 239476
rect 454404 239474 455004 239476
rect 490404 239474 491004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588080 239474 588680 239476
rect -2916 236476 -2316 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 198804 236476 199404 236478
rect 234804 236476 235404 236478
rect 270804 236476 271404 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586240 236476 586840 236478
rect -2916 236454 586840 236476
rect -2916 236218 -2734 236454
rect -2498 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 198986 236454
rect 199222 236218 234986 236454
rect 235222 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586422 236454
rect 586658 236218 586840 236454
rect -2916 236134 586840 236218
rect -2916 235898 -2734 236134
rect -2498 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 198986 236134
rect 199222 235898 234986 236134
rect 235222 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586422 236134
rect 586658 235898 586840 236134
rect -2916 235876 586840 235898
rect -2916 235874 -2316 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 198804 235874 199404 235876
rect 234804 235874 235404 235876
rect 270804 235874 271404 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586240 235874 586840 235876
rect -7516 229276 -6916 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 83604 229276 84204 229278
rect 119604 229276 120204 229278
rect 155604 229276 156204 229278
rect 191604 229276 192204 229278
rect 227604 229276 228204 229278
rect 263604 229276 264204 229278
rect 299604 229276 300204 229278
rect 335604 229276 336204 229278
rect 371604 229276 372204 229278
rect 407604 229276 408204 229278
rect 443604 229276 444204 229278
rect 479604 229276 480204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590840 229276 591440 229278
rect -8436 229254 592360 229276
rect -8436 229018 -7334 229254
rect -7098 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 83786 229254
rect 84022 229018 119786 229254
rect 120022 229018 155786 229254
rect 156022 229018 191786 229254
rect 192022 229018 227786 229254
rect 228022 229018 263786 229254
rect 264022 229018 299786 229254
rect 300022 229018 335786 229254
rect 336022 229018 371786 229254
rect 372022 229018 407786 229254
rect 408022 229018 443786 229254
rect 444022 229018 479786 229254
rect 480022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591022 229254
rect 591258 229018 592360 229254
rect -8436 228934 592360 229018
rect -8436 228698 -7334 228934
rect -7098 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 83786 228934
rect 84022 228698 119786 228934
rect 120022 228698 155786 228934
rect 156022 228698 191786 228934
rect 192022 228698 227786 228934
rect 228022 228698 263786 228934
rect 264022 228698 299786 228934
rect 300022 228698 335786 228934
rect 336022 228698 371786 228934
rect 372022 228698 407786 228934
rect 408022 228698 443786 228934
rect 444022 228698 479786 228934
rect 480022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591022 228934
rect 591258 228698 592360 228934
rect -8436 228676 592360 228698
rect -7516 228674 -6916 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 83604 228674 84204 228676
rect 119604 228674 120204 228676
rect 155604 228674 156204 228676
rect 191604 228674 192204 228676
rect 227604 228674 228204 228676
rect 263604 228674 264204 228676
rect 299604 228674 300204 228676
rect 335604 228674 336204 228676
rect 371604 228674 372204 228676
rect 407604 228674 408204 228676
rect 443604 228674 444204 228676
rect 479604 228674 480204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590840 228674 591440 228676
rect -5676 225676 -5076 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 116004 225676 116604 225678
rect 152004 225676 152604 225678
rect 188004 225676 188604 225678
rect 224004 225676 224604 225678
rect 260004 225676 260604 225678
rect 296004 225676 296604 225678
rect 332004 225676 332604 225678
rect 368004 225676 368604 225678
rect 404004 225676 404604 225678
rect 440004 225676 440604 225678
rect 476004 225676 476604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589000 225676 589600 225678
rect -6596 225654 590520 225676
rect -6596 225418 -5494 225654
rect -5258 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 116186 225654
rect 116422 225418 152186 225654
rect 152422 225418 188186 225654
rect 188422 225418 224186 225654
rect 224422 225418 260186 225654
rect 260422 225418 296186 225654
rect 296422 225418 332186 225654
rect 332422 225418 368186 225654
rect 368422 225418 404186 225654
rect 404422 225418 440186 225654
rect 440422 225418 476186 225654
rect 476422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589182 225654
rect 589418 225418 590520 225654
rect -6596 225334 590520 225418
rect -6596 225098 -5494 225334
rect -5258 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 116186 225334
rect 116422 225098 152186 225334
rect 152422 225098 188186 225334
rect 188422 225098 224186 225334
rect 224422 225098 260186 225334
rect 260422 225098 296186 225334
rect 296422 225098 332186 225334
rect 332422 225098 368186 225334
rect 368422 225098 404186 225334
rect 404422 225098 440186 225334
rect 440422 225098 476186 225334
rect 476422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589182 225334
rect 589418 225098 590520 225334
rect -6596 225076 590520 225098
rect -5676 225074 -5076 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 116004 225074 116604 225076
rect 152004 225074 152604 225076
rect 188004 225074 188604 225076
rect 224004 225074 224604 225076
rect 260004 225074 260604 225076
rect 296004 225074 296604 225076
rect 332004 225074 332604 225076
rect 368004 225074 368604 225076
rect 404004 225074 404604 225076
rect 440004 225074 440604 225076
rect 476004 225074 476604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589000 225074 589600 225076
rect -3836 222076 -3236 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 148404 222076 149004 222078
rect 184404 222076 185004 222078
rect 220404 222076 221004 222078
rect 256404 222076 257004 222078
rect 292404 222076 293004 222078
rect 328404 222076 329004 222078
rect 364404 222076 365004 222078
rect 400404 222076 401004 222078
rect 436404 222076 437004 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587160 222076 587760 222078
rect -4756 222054 588680 222076
rect -4756 221818 -3654 222054
rect -3418 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 148586 222054
rect 148822 221818 184586 222054
rect 184822 221818 220586 222054
rect 220822 221818 256586 222054
rect 256822 221818 292586 222054
rect 292822 221818 328586 222054
rect 328822 221818 364586 222054
rect 364822 221818 400586 222054
rect 400822 221818 436586 222054
rect 436822 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587342 222054
rect 587578 221818 588680 222054
rect -4756 221734 588680 221818
rect -4756 221498 -3654 221734
rect -3418 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 148586 221734
rect 148822 221498 184586 221734
rect 184822 221498 220586 221734
rect 220822 221498 256586 221734
rect 256822 221498 292586 221734
rect 292822 221498 328586 221734
rect 328822 221498 364586 221734
rect 364822 221498 400586 221734
rect 400822 221498 436586 221734
rect 436822 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587342 221734
rect 587578 221498 588680 221734
rect -4756 221476 588680 221498
rect -3836 221474 -3236 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 148404 221474 149004 221476
rect 184404 221474 185004 221476
rect 220404 221474 221004 221476
rect 256404 221474 257004 221476
rect 292404 221474 293004 221476
rect 328404 221474 329004 221476
rect 364404 221474 365004 221476
rect 400404 221474 401004 221476
rect 436404 221474 437004 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587160 221474 587760 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 144804 218476 145404 218478
rect 180804 218476 181404 218478
rect 216804 218476 217404 218478
rect 252804 218476 253404 218478
rect 288804 218476 289404 218478
rect 324804 218476 325404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2916 218454 586840 218476
rect -2916 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 180986 218454
rect 181222 218218 216986 218454
rect 217222 218218 252986 218454
rect 253222 218218 288986 218454
rect 289222 218218 324986 218454
rect 325222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586840 218454
rect -2916 218134 586840 218218
rect -2916 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 180986 218134
rect 181222 217898 216986 218134
rect 217222 217898 252986 218134
rect 253222 217898 288986 218134
rect 289222 217898 324986 218134
rect 325222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586840 218134
rect -2916 217876 586840 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 144804 217874 145404 217876
rect 180804 217874 181404 217876
rect 216804 217874 217404 217876
rect 252804 217874 253404 217876
rect 288804 217874 289404 217876
rect 324804 217874 325404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8436 211276 -7836 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 101604 211276 102204 211278
rect 137604 211276 138204 211278
rect 173604 211276 174204 211278
rect 209604 211276 210204 211278
rect 245604 211276 246204 211278
rect 281604 211276 282204 211278
rect 317604 211276 318204 211278
rect 353604 211276 354204 211278
rect 389604 211276 390204 211278
rect 425604 211276 426204 211278
rect 461604 211276 462204 211278
rect 497604 211276 498204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591760 211276 592360 211278
rect -8436 211254 592360 211276
rect -8436 211018 -8254 211254
rect -8018 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 101786 211254
rect 102022 211018 137786 211254
rect 138022 211018 173786 211254
rect 174022 211018 209786 211254
rect 210022 211018 245786 211254
rect 246022 211018 281786 211254
rect 282022 211018 317786 211254
rect 318022 211018 353786 211254
rect 354022 211018 389786 211254
rect 390022 211018 425786 211254
rect 426022 211018 461786 211254
rect 462022 211018 497786 211254
rect 498022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 591942 211254
rect 592178 211018 592360 211254
rect -8436 210934 592360 211018
rect -8436 210698 -8254 210934
rect -8018 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 101786 210934
rect 102022 210698 137786 210934
rect 138022 210698 173786 210934
rect 174022 210698 209786 210934
rect 210022 210698 245786 210934
rect 246022 210698 281786 210934
rect 282022 210698 317786 210934
rect 318022 210698 353786 210934
rect 354022 210698 389786 210934
rect 390022 210698 425786 210934
rect 426022 210698 461786 210934
rect 462022 210698 497786 210934
rect 498022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 591942 210934
rect 592178 210698 592360 210934
rect -8436 210676 592360 210698
rect -8436 210674 -7836 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 101604 210674 102204 210676
rect 137604 210674 138204 210676
rect 173604 210674 174204 210676
rect 209604 210674 210204 210676
rect 245604 210674 246204 210676
rect 281604 210674 282204 210676
rect 317604 210674 318204 210676
rect 353604 210674 354204 210676
rect 389604 210674 390204 210676
rect 425604 210674 426204 210676
rect 461604 210674 462204 210676
rect 497604 210674 498204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591760 210674 592360 210676
rect -6596 207676 -5996 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 98004 207676 98604 207678
rect 134004 207676 134604 207678
rect 170004 207676 170604 207678
rect 206004 207676 206604 207678
rect 242004 207676 242604 207678
rect 278004 207676 278604 207678
rect 314004 207676 314604 207678
rect 350004 207676 350604 207678
rect 386004 207676 386604 207678
rect 422004 207676 422604 207678
rect 458004 207676 458604 207678
rect 494004 207676 494604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 589920 207676 590520 207678
rect -6596 207654 590520 207676
rect -6596 207418 -6414 207654
rect -6178 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 98186 207654
rect 98422 207418 134186 207654
rect 134422 207418 170186 207654
rect 170422 207418 206186 207654
rect 206422 207418 242186 207654
rect 242422 207418 278186 207654
rect 278422 207418 314186 207654
rect 314422 207418 350186 207654
rect 350422 207418 386186 207654
rect 386422 207418 422186 207654
rect 422422 207418 458186 207654
rect 458422 207418 494186 207654
rect 494422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590102 207654
rect 590338 207418 590520 207654
rect -6596 207334 590520 207418
rect -6596 207098 -6414 207334
rect -6178 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 98186 207334
rect 98422 207098 134186 207334
rect 134422 207098 170186 207334
rect 170422 207098 206186 207334
rect 206422 207098 242186 207334
rect 242422 207098 278186 207334
rect 278422 207098 314186 207334
rect 314422 207098 350186 207334
rect 350422 207098 386186 207334
rect 386422 207098 422186 207334
rect 422422 207098 458186 207334
rect 458422 207098 494186 207334
rect 494422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590102 207334
rect 590338 207098 590520 207334
rect -6596 207076 590520 207098
rect -6596 207074 -5996 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 98004 207074 98604 207076
rect 134004 207074 134604 207076
rect 170004 207074 170604 207076
rect 206004 207074 206604 207076
rect 242004 207074 242604 207076
rect 278004 207074 278604 207076
rect 314004 207074 314604 207076
rect 350004 207074 350604 207076
rect 386004 207074 386604 207076
rect 422004 207074 422604 207076
rect 458004 207074 458604 207076
rect 494004 207074 494604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 589920 207074 590520 207076
rect -4756 204076 -4156 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 166404 204076 167004 204078
rect 202404 204076 203004 204078
rect 238404 204076 239004 204078
rect 274404 204076 275004 204078
rect 310404 204076 311004 204078
rect 346404 204076 347004 204078
rect 382404 204076 383004 204078
rect 418404 204076 419004 204078
rect 454404 204076 455004 204078
rect 490404 204076 491004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588080 204076 588680 204078
rect -4756 204054 588680 204076
rect -4756 203818 -4574 204054
rect -4338 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 166586 204054
rect 166822 203818 202586 204054
rect 202822 203818 238586 204054
rect 238822 203818 274586 204054
rect 274822 203818 310586 204054
rect 310822 203818 346586 204054
rect 346822 203818 382586 204054
rect 382822 203818 418586 204054
rect 418822 203818 454586 204054
rect 454822 203818 490586 204054
rect 490822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588262 204054
rect 588498 203818 588680 204054
rect -4756 203734 588680 203818
rect -4756 203498 -4574 203734
rect -4338 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 166586 203734
rect 166822 203498 202586 203734
rect 202822 203498 238586 203734
rect 238822 203498 274586 203734
rect 274822 203498 310586 203734
rect 310822 203498 346586 203734
rect 346822 203498 382586 203734
rect 382822 203498 418586 203734
rect 418822 203498 454586 203734
rect 454822 203498 490586 203734
rect 490822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588262 203734
rect 588498 203498 588680 203734
rect -4756 203476 588680 203498
rect -4756 203474 -4156 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 166404 203474 167004 203476
rect 202404 203474 203004 203476
rect 238404 203474 239004 203476
rect 274404 203474 275004 203476
rect 310404 203474 311004 203476
rect 346404 203474 347004 203476
rect 382404 203474 383004 203476
rect 418404 203474 419004 203476
rect 454404 203474 455004 203476
rect 490404 203474 491004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588080 203474 588680 203476
rect -2916 200476 -2316 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 162804 200476 163404 200478
rect 198804 200476 199404 200478
rect 234804 200476 235404 200478
rect 270804 200476 271404 200478
rect 306804 200476 307404 200478
rect 342804 200476 343404 200478
rect 378804 200476 379404 200478
rect 414804 200476 415404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586240 200476 586840 200478
rect -2916 200454 586840 200476
rect -2916 200218 -2734 200454
rect -2498 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 162986 200454
rect 163222 200218 198986 200454
rect 199222 200218 234986 200454
rect 235222 200218 270986 200454
rect 271222 200218 306986 200454
rect 307222 200218 342986 200454
rect 343222 200218 378986 200454
rect 379222 200218 414986 200454
rect 415222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586422 200454
rect 586658 200218 586840 200454
rect -2916 200134 586840 200218
rect -2916 199898 -2734 200134
rect -2498 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 162986 200134
rect 163222 199898 198986 200134
rect 199222 199898 234986 200134
rect 235222 199898 270986 200134
rect 271222 199898 306986 200134
rect 307222 199898 342986 200134
rect 343222 199898 378986 200134
rect 379222 199898 414986 200134
rect 415222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586422 200134
rect 586658 199898 586840 200134
rect -2916 199876 586840 199898
rect -2916 199874 -2316 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 162804 199874 163404 199876
rect 198804 199874 199404 199876
rect 234804 199874 235404 199876
rect 270804 199874 271404 199876
rect 306804 199874 307404 199876
rect 342804 199874 343404 199876
rect 378804 199874 379404 199876
rect 414804 199874 415404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586240 199874 586840 199876
rect -7516 193276 -6916 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 155604 193276 156204 193278
rect 191604 193276 192204 193278
rect 227604 193276 228204 193278
rect 263604 193276 264204 193278
rect 299604 193276 300204 193278
rect 335604 193276 336204 193278
rect 371604 193276 372204 193278
rect 407604 193276 408204 193278
rect 443604 193276 444204 193278
rect 479604 193276 480204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590840 193276 591440 193278
rect -8436 193254 592360 193276
rect -8436 193018 -7334 193254
rect -7098 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 155786 193254
rect 156022 193018 191786 193254
rect 192022 193018 227786 193254
rect 228022 193018 263786 193254
rect 264022 193018 299786 193254
rect 300022 193018 335786 193254
rect 336022 193018 371786 193254
rect 372022 193018 407786 193254
rect 408022 193018 443786 193254
rect 444022 193018 479786 193254
rect 480022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591022 193254
rect 591258 193018 592360 193254
rect -8436 192934 592360 193018
rect -8436 192698 -7334 192934
rect -7098 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 155786 192934
rect 156022 192698 191786 192934
rect 192022 192698 227786 192934
rect 228022 192698 263786 192934
rect 264022 192698 299786 192934
rect 300022 192698 335786 192934
rect 336022 192698 371786 192934
rect 372022 192698 407786 192934
rect 408022 192698 443786 192934
rect 444022 192698 479786 192934
rect 480022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591022 192934
rect 591258 192698 592360 192934
rect -8436 192676 592360 192698
rect -7516 192674 -6916 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 155604 192674 156204 192676
rect 191604 192674 192204 192676
rect 227604 192674 228204 192676
rect 263604 192674 264204 192676
rect 299604 192674 300204 192676
rect 335604 192674 336204 192676
rect 371604 192674 372204 192676
rect 407604 192674 408204 192676
rect 443604 192674 444204 192676
rect 479604 192674 480204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590840 192674 591440 192676
rect -5676 189676 -5076 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 152004 189676 152604 189678
rect 188004 189676 188604 189678
rect 224004 189676 224604 189678
rect 260004 189676 260604 189678
rect 296004 189676 296604 189678
rect 332004 189676 332604 189678
rect 368004 189676 368604 189678
rect 404004 189676 404604 189678
rect 440004 189676 440604 189678
rect 476004 189676 476604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589000 189676 589600 189678
rect -6596 189654 590520 189676
rect -6596 189418 -5494 189654
rect -5258 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 152186 189654
rect 152422 189418 188186 189654
rect 188422 189418 224186 189654
rect 224422 189418 260186 189654
rect 260422 189418 296186 189654
rect 296422 189418 332186 189654
rect 332422 189418 368186 189654
rect 368422 189418 404186 189654
rect 404422 189418 440186 189654
rect 440422 189418 476186 189654
rect 476422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589182 189654
rect 589418 189418 590520 189654
rect -6596 189334 590520 189418
rect -6596 189098 -5494 189334
rect -5258 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 152186 189334
rect 152422 189098 188186 189334
rect 188422 189098 224186 189334
rect 224422 189098 260186 189334
rect 260422 189098 296186 189334
rect 296422 189098 332186 189334
rect 332422 189098 368186 189334
rect 368422 189098 404186 189334
rect 404422 189098 440186 189334
rect 440422 189098 476186 189334
rect 476422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589182 189334
rect 589418 189098 590520 189334
rect -6596 189076 590520 189098
rect -5676 189074 -5076 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 152004 189074 152604 189076
rect 188004 189074 188604 189076
rect 224004 189074 224604 189076
rect 260004 189074 260604 189076
rect 296004 189074 296604 189076
rect 332004 189074 332604 189076
rect 368004 189074 368604 189076
rect 404004 189074 404604 189076
rect 440004 189074 440604 189076
rect 476004 189074 476604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589000 189074 589600 189076
rect -3836 186076 -3236 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 148404 186076 149004 186078
rect 184404 186076 185004 186078
rect 220404 186076 221004 186078
rect 256404 186076 257004 186078
rect 292404 186076 293004 186078
rect 328404 186076 329004 186078
rect 364404 186076 365004 186078
rect 400404 186076 401004 186078
rect 436404 186076 437004 186078
rect 472404 186076 473004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587160 186076 587760 186078
rect -4756 186054 588680 186076
rect -4756 185818 -3654 186054
rect -3418 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 148586 186054
rect 148822 185818 184586 186054
rect 184822 185818 220586 186054
rect 220822 185818 256586 186054
rect 256822 185818 292586 186054
rect 292822 185818 328586 186054
rect 328822 185818 364586 186054
rect 364822 185818 400586 186054
rect 400822 185818 436586 186054
rect 436822 185818 472586 186054
rect 472822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587342 186054
rect 587578 185818 588680 186054
rect -4756 185734 588680 185818
rect -4756 185498 -3654 185734
rect -3418 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 148586 185734
rect 148822 185498 184586 185734
rect 184822 185498 220586 185734
rect 220822 185498 256586 185734
rect 256822 185498 292586 185734
rect 292822 185498 328586 185734
rect 328822 185498 364586 185734
rect 364822 185498 400586 185734
rect 400822 185498 436586 185734
rect 436822 185498 472586 185734
rect 472822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587342 185734
rect 587578 185498 588680 185734
rect -4756 185476 588680 185498
rect -3836 185474 -3236 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 148404 185474 149004 185476
rect 184404 185474 185004 185476
rect 220404 185474 221004 185476
rect 256404 185474 257004 185476
rect 292404 185474 293004 185476
rect 328404 185474 329004 185476
rect 364404 185474 365004 185476
rect 400404 185474 401004 185476
rect 436404 185474 437004 185476
rect 472404 185474 473004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587160 185474 587760 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 180804 182476 181404 182478
rect 216804 182476 217404 182478
rect 252804 182476 253404 182478
rect 288804 182476 289404 182478
rect 324804 182476 325404 182478
rect 360804 182476 361404 182478
rect 396804 182476 397404 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2916 182454 586840 182476
rect -2916 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 324986 182454
rect 325222 182218 360986 182454
rect 361222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586840 182454
rect -2916 182134 586840 182218
rect -2916 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 324986 182134
rect 325222 181898 360986 182134
rect 361222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586840 182134
rect -2916 181876 586840 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 180804 181874 181404 181876
rect 216804 181874 217404 181876
rect 252804 181874 253404 181876
rect 288804 181874 289404 181876
rect 324804 181874 325404 181876
rect 360804 181874 361404 181876
rect 396804 181874 397404 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8436 175276 -7836 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 137604 175276 138204 175278
rect 173604 175276 174204 175278
rect 209604 175276 210204 175278
rect 245604 175276 246204 175278
rect 281604 175276 282204 175278
rect 317604 175276 318204 175278
rect 353604 175276 354204 175278
rect 389604 175276 390204 175278
rect 425604 175276 426204 175278
rect 461604 175276 462204 175278
rect 497604 175276 498204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591760 175276 592360 175278
rect -8436 175254 592360 175276
rect -8436 175018 -8254 175254
rect -8018 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 137786 175254
rect 138022 175018 173786 175254
rect 174022 175018 209786 175254
rect 210022 175018 245786 175254
rect 246022 175018 281786 175254
rect 282022 175018 317786 175254
rect 318022 175018 353786 175254
rect 354022 175018 389786 175254
rect 390022 175018 425786 175254
rect 426022 175018 461786 175254
rect 462022 175018 497786 175254
rect 498022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 591942 175254
rect 592178 175018 592360 175254
rect -8436 174934 592360 175018
rect -8436 174698 -8254 174934
rect -8018 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 137786 174934
rect 138022 174698 173786 174934
rect 174022 174698 209786 174934
rect 210022 174698 245786 174934
rect 246022 174698 281786 174934
rect 282022 174698 317786 174934
rect 318022 174698 353786 174934
rect 354022 174698 389786 174934
rect 390022 174698 425786 174934
rect 426022 174698 461786 174934
rect 462022 174698 497786 174934
rect 498022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 591942 174934
rect 592178 174698 592360 174934
rect -8436 174676 592360 174698
rect -8436 174674 -7836 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 137604 174674 138204 174676
rect 173604 174674 174204 174676
rect 209604 174674 210204 174676
rect 245604 174674 246204 174676
rect 281604 174674 282204 174676
rect 317604 174674 318204 174676
rect 353604 174674 354204 174676
rect 389604 174674 390204 174676
rect 425604 174674 426204 174676
rect 461604 174674 462204 174676
rect 497604 174674 498204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591760 174674 592360 174676
rect -6596 171676 -5996 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 134004 171676 134604 171678
rect 170004 171676 170604 171678
rect 206004 171676 206604 171678
rect 242004 171676 242604 171678
rect 278004 171676 278604 171678
rect 314004 171676 314604 171678
rect 350004 171676 350604 171678
rect 386004 171676 386604 171678
rect 422004 171676 422604 171678
rect 458004 171676 458604 171678
rect 494004 171676 494604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 589920 171676 590520 171678
rect -6596 171654 590520 171676
rect -6596 171418 -6414 171654
rect -6178 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 134186 171654
rect 134422 171418 170186 171654
rect 170422 171418 206186 171654
rect 206422 171418 242186 171654
rect 242422 171418 278186 171654
rect 278422 171418 314186 171654
rect 314422 171418 350186 171654
rect 350422 171418 386186 171654
rect 386422 171418 422186 171654
rect 422422 171418 458186 171654
rect 458422 171418 494186 171654
rect 494422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590102 171654
rect 590338 171418 590520 171654
rect -6596 171334 590520 171418
rect -6596 171098 -6414 171334
rect -6178 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 134186 171334
rect 134422 171098 170186 171334
rect 170422 171098 206186 171334
rect 206422 171098 242186 171334
rect 242422 171098 278186 171334
rect 278422 171098 314186 171334
rect 314422 171098 350186 171334
rect 350422 171098 386186 171334
rect 386422 171098 422186 171334
rect 422422 171098 458186 171334
rect 458422 171098 494186 171334
rect 494422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590102 171334
rect 590338 171098 590520 171334
rect -6596 171076 590520 171098
rect -6596 171074 -5996 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 134004 171074 134604 171076
rect 170004 171074 170604 171076
rect 206004 171074 206604 171076
rect 242004 171074 242604 171076
rect 278004 171074 278604 171076
rect 314004 171074 314604 171076
rect 350004 171074 350604 171076
rect 386004 171074 386604 171076
rect 422004 171074 422604 171076
rect 458004 171074 458604 171076
rect 494004 171074 494604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 589920 171074 590520 171076
rect -4756 168076 -4156 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 166404 168076 167004 168078
rect 202404 168076 203004 168078
rect 238404 168076 239004 168078
rect 274404 168076 275004 168078
rect 310404 168076 311004 168078
rect 346404 168076 347004 168078
rect 382404 168076 383004 168078
rect 418404 168076 419004 168078
rect 454404 168076 455004 168078
rect 490404 168076 491004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588080 168076 588680 168078
rect -4756 168054 588680 168076
rect -4756 167818 -4574 168054
rect -4338 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 166586 168054
rect 166822 167818 202586 168054
rect 202822 167818 238586 168054
rect 238822 167818 274586 168054
rect 274822 167818 310586 168054
rect 310822 167818 346586 168054
rect 346822 167818 382586 168054
rect 382822 167818 418586 168054
rect 418822 167818 454586 168054
rect 454822 167818 490586 168054
rect 490822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588262 168054
rect 588498 167818 588680 168054
rect -4756 167734 588680 167818
rect -4756 167498 -4574 167734
rect -4338 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 166586 167734
rect 166822 167498 202586 167734
rect 202822 167498 238586 167734
rect 238822 167498 274586 167734
rect 274822 167498 310586 167734
rect 310822 167498 346586 167734
rect 346822 167498 382586 167734
rect 382822 167498 418586 167734
rect 418822 167498 454586 167734
rect 454822 167498 490586 167734
rect 490822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588262 167734
rect 588498 167498 588680 167734
rect -4756 167476 588680 167498
rect -4756 167474 -4156 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 166404 167474 167004 167476
rect 202404 167474 203004 167476
rect 238404 167474 239004 167476
rect 274404 167474 275004 167476
rect 310404 167474 311004 167476
rect 346404 167474 347004 167476
rect 382404 167474 383004 167476
rect 418404 167474 419004 167476
rect 454404 167474 455004 167476
rect 490404 167474 491004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588080 167474 588680 167476
rect -2916 164476 -2316 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 342804 164476 343404 164478
rect 378804 164476 379404 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586240 164476 586840 164478
rect -2916 164454 586840 164476
rect -2916 164218 -2734 164454
rect -2498 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586422 164454
rect 586658 164218 586840 164454
rect -2916 164134 586840 164218
rect -2916 163898 -2734 164134
rect -2498 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586422 164134
rect 586658 163898 586840 164134
rect -2916 163876 586840 163898
rect -2916 163874 -2316 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 342804 163874 343404 163876
rect 378804 163874 379404 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586240 163874 586840 163876
rect -7516 157276 -6916 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 155604 157276 156204 157278
rect 191604 157276 192204 157278
rect 227604 157276 228204 157278
rect 263604 157276 264204 157278
rect 299604 157276 300204 157278
rect 335604 157276 336204 157278
rect 371604 157276 372204 157278
rect 407604 157276 408204 157278
rect 443604 157276 444204 157278
rect 479604 157276 480204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590840 157276 591440 157278
rect -8436 157254 592360 157276
rect -8436 157018 -7334 157254
rect -7098 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 155786 157254
rect 156022 157018 191786 157254
rect 192022 157018 227786 157254
rect 228022 157018 263786 157254
rect 264022 157018 299786 157254
rect 300022 157018 335786 157254
rect 336022 157018 371786 157254
rect 372022 157018 407786 157254
rect 408022 157018 443786 157254
rect 444022 157018 479786 157254
rect 480022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591022 157254
rect 591258 157018 592360 157254
rect -8436 156934 592360 157018
rect -8436 156698 -7334 156934
rect -7098 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 155786 156934
rect 156022 156698 191786 156934
rect 192022 156698 227786 156934
rect 228022 156698 263786 156934
rect 264022 156698 299786 156934
rect 300022 156698 335786 156934
rect 336022 156698 371786 156934
rect 372022 156698 407786 156934
rect 408022 156698 443786 156934
rect 444022 156698 479786 156934
rect 480022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591022 156934
rect 591258 156698 592360 156934
rect -8436 156676 592360 156698
rect -7516 156674 -6916 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 155604 156674 156204 156676
rect 191604 156674 192204 156676
rect 227604 156674 228204 156676
rect 263604 156674 264204 156676
rect 299604 156674 300204 156676
rect 335604 156674 336204 156676
rect 371604 156674 372204 156676
rect 407604 156674 408204 156676
rect 443604 156674 444204 156676
rect 479604 156674 480204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590840 156674 591440 156676
rect -5676 153676 -5076 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 152004 153676 152604 153678
rect 188004 153676 188604 153678
rect 224004 153676 224604 153678
rect 260004 153676 260604 153678
rect 296004 153676 296604 153678
rect 332004 153676 332604 153678
rect 368004 153676 368604 153678
rect 404004 153676 404604 153678
rect 440004 153676 440604 153678
rect 476004 153676 476604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589000 153676 589600 153678
rect -6596 153654 590520 153676
rect -6596 153418 -5494 153654
rect -5258 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 152186 153654
rect 152422 153418 188186 153654
rect 188422 153418 224186 153654
rect 224422 153418 260186 153654
rect 260422 153418 296186 153654
rect 296422 153418 332186 153654
rect 332422 153418 368186 153654
rect 368422 153418 404186 153654
rect 404422 153418 440186 153654
rect 440422 153418 476186 153654
rect 476422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589182 153654
rect 589418 153418 590520 153654
rect -6596 153334 590520 153418
rect -6596 153098 -5494 153334
rect -5258 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 152186 153334
rect 152422 153098 188186 153334
rect 188422 153098 224186 153334
rect 224422 153098 260186 153334
rect 260422 153098 296186 153334
rect 296422 153098 332186 153334
rect 332422 153098 368186 153334
rect 368422 153098 404186 153334
rect 404422 153098 440186 153334
rect 440422 153098 476186 153334
rect 476422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589182 153334
rect 589418 153098 590520 153334
rect -6596 153076 590520 153098
rect -5676 153074 -5076 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 152004 153074 152604 153076
rect 188004 153074 188604 153076
rect 224004 153074 224604 153076
rect 260004 153074 260604 153076
rect 296004 153074 296604 153076
rect 332004 153074 332604 153076
rect 368004 153074 368604 153076
rect 404004 153074 404604 153076
rect 440004 153074 440604 153076
rect 476004 153074 476604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589000 153074 589600 153076
rect -3836 150076 -3236 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 148404 150076 149004 150078
rect 184404 150076 185004 150078
rect 220404 150076 221004 150078
rect 256404 150076 257004 150078
rect 292404 150076 293004 150078
rect 328404 150076 329004 150078
rect 364404 150076 365004 150078
rect 400404 150076 401004 150078
rect 436404 150076 437004 150078
rect 472404 150076 473004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587160 150076 587760 150078
rect -4756 150054 588680 150076
rect -4756 149818 -3654 150054
rect -3418 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 148586 150054
rect 148822 149818 184586 150054
rect 184822 149818 220586 150054
rect 220822 149818 256586 150054
rect 256822 149818 292586 150054
rect 292822 149818 328586 150054
rect 328822 149818 364586 150054
rect 364822 149818 400586 150054
rect 400822 149818 436586 150054
rect 436822 149818 472586 150054
rect 472822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587342 150054
rect 587578 149818 588680 150054
rect -4756 149734 588680 149818
rect -4756 149498 -3654 149734
rect -3418 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 148586 149734
rect 148822 149498 184586 149734
rect 184822 149498 220586 149734
rect 220822 149498 256586 149734
rect 256822 149498 292586 149734
rect 292822 149498 328586 149734
rect 328822 149498 364586 149734
rect 364822 149498 400586 149734
rect 400822 149498 436586 149734
rect 436822 149498 472586 149734
rect 472822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587342 149734
rect 587578 149498 588680 149734
rect -4756 149476 588680 149498
rect -3836 149474 -3236 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 148404 149474 149004 149476
rect 184404 149474 185004 149476
rect 220404 149474 221004 149476
rect 256404 149474 257004 149476
rect 292404 149474 293004 149476
rect 328404 149474 329004 149476
rect 364404 149474 365004 149476
rect 400404 149474 401004 149476
rect 436404 149474 437004 149476
rect 472404 149474 473004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587160 149474 587760 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 324804 146476 325404 146478
rect 360804 146476 361404 146478
rect 396804 146476 397404 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2916 146454 586840 146476
rect -2916 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 324986 146454
rect 325222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586840 146454
rect -2916 146134 586840 146218
rect -2916 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 324986 146134
rect 325222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586840 146134
rect -2916 145876 586840 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 324804 145874 325404 145876
rect 360804 145874 361404 145876
rect 396804 145874 397404 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8436 139276 -7836 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 137604 139276 138204 139278
rect 173604 139276 174204 139278
rect 209604 139276 210204 139278
rect 245604 139276 246204 139278
rect 281604 139276 282204 139278
rect 317604 139276 318204 139278
rect 353604 139276 354204 139278
rect 389604 139276 390204 139278
rect 425604 139276 426204 139278
rect 461604 139276 462204 139278
rect 497604 139276 498204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591760 139276 592360 139278
rect -8436 139254 592360 139276
rect -8436 139018 -8254 139254
rect -8018 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 137786 139254
rect 138022 139018 173786 139254
rect 174022 139018 209786 139254
rect 210022 139018 245786 139254
rect 246022 139018 281786 139254
rect 282022 139018 317786 139254
rect 318022 139018 353786 139254
rect 354022 139018 389786 139254
rect 390022 139018 425786 139254
rect 426022 139018 461786 139254
rect 462022 139018 497786 139254
rect 498022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 591942 139254
rect 592178 139018 592360 139254
rect -8436 138934 592360 139018
rect -8436 138698 -8254 138934
rect -8018 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 137786 138934
rect 138022 138698 173786 138934
rect 174022 138698 209786 138934
rect 210022 138698 245786 138934
rect 246022 138698 281786 138934
rect 282022 138698 317786 138934
rect 318022 138698 353786 138934
rect 354022 138698 389786 138934
rect 390022 138698 425786 138934
rect 426022 138698 461786 138934
rect 462022 138698 497786 138934
rect 498022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 591942 138934
rect 592178 138698 592360 138934
rect -8436 138676 592360 138698
rect -8436 138674 -7836 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 137604 138674 138204 138676
rect 173604 138674 174204 138676
rect 209604 138674 210204 138676
rect 245604 138674 246204 138676
rect 281604 138674 282204 138676
rect 317604 138674 318204 138676
rect 353604 138674 354204 138676
rect 389604 138674 390204 138676
rect 425604 138674 426204 138676
rect 461604 138674 462204 138676
rect 497604 138674 498204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591760 138674 592360 138676
rect -6596 135676 -5996 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 134004 135676 134604 135678
rect 170004 135676 170604 135678
rect 206004 135676 206604 135678
rect 242004 135676 242604 135678
rect 278004 135676 278604 135678
rect 314004 135676 314604 135678
rect 350004 135676 350604 135678
rect 386004 135676 386604 135678
rect 422004 135676 422604 135678
rect 458004 135676 458604 135678
rect 494004 135676 494604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 589920 135676 590520 135678
rect -6596 135654 590520 135676
rect -6596 135418 -6414 135654
rect -6178 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 134186 135654
rect 134422 135418 170186 135654
rect 170422 135418 206186 135654
rect 206422 135418 242186 135654
rect 242422 135418 278186 135654
rect 278422 135418 314186 135654
rect 314422 135418 350186 135654
rect 350422 135418 386186 135654
rect 386422 135418 422186 135654
rect 422422 135418 458186 135654
rect 458422 135418 494186 135654
rect 494422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590102 135654
rect 590338 135418 590520 135654
rect -6596 135334 590520 135418
rect -6596 135098 -6414 135334
rect -6178 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 134186 135334
rect 134422 135098 170186 135334
rect 170422 135098 206186 135334
rect 206422 135098 242186 135334
rect 242422 135098 278186 135334
rect 278422 135098 314186 135334
rect 314422 135098 350186 135334
rect 350422 135098 386186 135334
rect 386422 135098 422186 135334
rect 422422 135098 458186 135334
rect 458422 135098 494186 135334
rect 494422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590102 135334
rect 590338 135098 590520 135334
rect -6596 135076 590520 135098
rect -6596 135074 -5996 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 134004 135074 134604 135076
rect 170004 135074 170604 135076
rect 206004 135074 206604 135076
rect 242004 135074 242604 135076
rect 278004 135074 278604 135076
rect 314004 135074 314604 135076
rect 350004 135074 350604 135076
rect 386004 135074 386604 135076
rect 422004 135074 422604 135076
rect 458004 135074 458604 135076
rect 494004 135074 494604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 589920 135074 590520 135076
rect -4756 132076 -4156 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 166404 132076 167004 132078
rect 202404 132076 203004 132078
rect 238404 132076 239004 132078
rect 274404 132076 275004 132078
rect 310404 132076 311004 132078
rect 346404 132076 347004 132078
rect 382404 132076 383004 132078
rect 418404 132076 419004 132078
rect 454404 132076 455004 132078
rect 490404 132076 491004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588080 132076 588680 132078
rect -4756 132054 588680 132076
rect -4756 131818 -4574 132054
rect -4338 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 166586 132054
rect 166822 131818 202586 132054
rect 202822 131818 238586 132054
rect 238822 131818 274586 132054
rect 274822 131818 310586 132054
rect 310822 131818 346586 132054
rect 346822 131818 382586 132054
rect 382822 131818 418586 132054
rect 418822 131818 454586 132054
rect 454822 131818 490586 132054
rect 490822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588262 132054
rect 588498 131818 588680 132054
rect -4756 131734 588680 131818
rect -4756 131498 -4574 131734
rect -4338 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 166586 131734
rect 166822 131498 202586 131734
rect 202822 131498 238586 131734
rect 238822 131498 274586 131734
rect 274822 131498 310586 131734
rect 310822 131498 346586 131734
rect 346822 131498 382586 131734
rect 382822 131498 418586 131734
rect 418822 131498 454586 131734
rect 454822 131498 490586 131734
rect 490822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588262 131734
rect 588498 131498 588680 131734
rect -4756 131476 588680 131498
rect -4756 131474 -4156 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 166404 131474 167004 131476
rect 202404 131474 203004 131476
rect 238404 131474 239004 131476
rect 274404 131474 275004 131476
rect 310404 131474 311004 131476
rect 346404 131474 347004 131476
rect 382404 131474 383004 131476
rect 418404 131474 419004 131476
rect 454404 131474 455004 131476
rect 490404 131474 491004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588080 131474 588680 131476
rect -2916 128476 -2316 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 306804 128476 307404 128478
rect 342804 128476 343404 128478
rect 378804 128476 379404 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586240 128476 586840 128478
rect -2916 128454 586840 128476
rect -2916 128218 -2734 128454
rect -2498 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586422 128454
rect 586658 128218 586840 128454
rect -2916 128134 586840 128218
rect -2916 127898 -2734 128134
rect -2498 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586422 128134
rect 586658 127898 586840 128134
rect -2916 127876 586840 127898
rect -2916 127874 -2316 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 306804 127874 307404 127876
rect 342804 127874 343404 127876
rect 378804 127874 379404 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586240 127874 586840 127876
rect -7516 121276 -6916 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 155604 121276 156204 121278
rect 191604 121276 192204 121278
rect 227604 121276 228204 121278
rect 263604 121276 264204 121278
rect 299604 121276 300204 121278
rect 335604 121276 336204 121278
rect 371604 121276 372204 121278
rect 407604 121276 408204 121278
rect 443604 121276 444204 121278
rect 479604 121276 480204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590840 121276 591440 121278
rect -8436 121254 592360 121276
rect -8436 121018 -7334 121254
rect -7098 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 155786 121254
rect 156022 121018 191786 121254
rect 192022 121018 227786 121254
rect 228022 121018 263786 121254
rect 264022 121018 299786 121254
rect 300022 121018 335786 121254
rect 336022 121018 371786 121254
rect 372022 121018 407786 121254
rect 408022 121018 443786 121254
rect 444022 121018 479786 121254
rect 480022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591022 121254
rect 591258 121018 592360 121254
rect -8436 120934 592360 121018
rect -8436 120698 -7334 120934
rect -7098 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 155786 120934
rect 156022 120698 191786 120934
rect 192022 120698 227786 120934
rect 228022 120698 263786 120934
rect 264022 120698 299786 120934
rect 300022 120698 335786 120934
rect 336022 120698 371786 120934
rect 372022 120698 407786 120934
rect 408022 120698 443786 120934
rect 444022 120698 479786 120934
rect 480022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591022 120934
rect 591258 120698 592360 120934
rect -8436 120676 592360 120698
rect -7516 120674 -6916 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 155604 120674 156204 120676
rect 191604 120674 192204 120676
rect 227604 120674 228204 120676
rect 263604 120674 264204 120676
rect 299604 120674 300204 120676
rect 335604 120674 336204 120676
rect 371604 120674 372204 120676
rect 407604 120674 408204 120676
rect 443604 120674 444204 120676
rect 479604 120674 480204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590840 120674 591440 120676
rect -5676 117676 -5076 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 332004 117676 332604 117678
rect 368004 117676 368604 117678
rect 404004 117676 404604 117678
rect 440004 117676 440604 117678
rect 476004 117676 476604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589000 117676 589600 117678
rect -6596 117654 590520 117676
rect -6596 117418 -5494 117654
rect -5258 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 332186 117654
rect 332422 117418 368186 117654
rect 368422 117418 404186 117654
rect 404422 117418 440186 117654
rect 440422 117418 476186 117654
rect 476422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589182 117654
rect 589418 117418 590520 117654
rect -6596 117334 590520 117418
rect -6596 117098 -5494 117334
rect -5258 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 332186 117334
rect 332422 117098 368186 117334
rect 368422 117098 404186 117334
rect 404422 117098 440186 117334
rect 440422 117098 476186 117334
rect 476422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589182 117334
rect 589418 117098 590520 117334
rect -6596 117076 590520 117098
rect -5676 117074 -5076 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 332004 117074 332604 117076
rect 368004 117074 368604 117076
rect 404004 117074 404604 117076
rect 440004 117074 440604 117076
rect 476004 117074 476604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589000 117074 589600 117076
rect -3836 114076 -3236 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 328404 114076 329004 114078
rect 364404 114076 365004 114078
rect 400404 114076 401004 114078
rect 436404 114076 437004 114078
rect 472404 114076 473004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587160 114076 587760 114078
rect -4756 114054 588680 114076
rect -4756 113818 -3654 114054
rect -3418 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 328586 114054
rect 328822 113818 364586 114054
rect 364822 113818 400586 114054
rect 400822 113818 436586 114054
rect 436822 113818 472586 114054
rect 472822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587342 114054
rect 587578 113818 588680 114054
rect -4756 113734 588680 113818
rect -4756 113498 -3654 113734
rect -3418 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 328586 113734
rect 328822 113498 364586 113734
rect 364822 113498 400586 113734
rect 400822 113498 436586 113734
rect 436822 113498 472586 113734
rect 472822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587342 113734
rect 587578 113498 588680 113734
rect -4756 113476 588680 113498
rect -3836 113474 -3236 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 328404 113474 329004 113476
rect 364404 113474 365004 113476
rect 400404 113474 401004 113476
rect 436404 113474 437004 113476
rect 472404 113474 473004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587160 113474 587760 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2916 110454 586840 110476
rect -2916 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586840 110454
rect -2916 110134 586840 110218
rect -2916 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586840 110134
rect -2916 109876 586840 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8436 103276 -7836 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 317604 103276 318204 103278
rect 353604 103276 354204 103278
rect 389604 103276 390204 103278
rect 425604 103276 426204 103278
rect 461604 103276 462204 103278
rect 497604 103276 498204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591760 103276 592360 103278
rect -8436 103254 592360 103276
rect -8436 103018 -8254 103254
rect -8018 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 317786 103254
rect 318022 103018 353786 103254
rect 354022 103018 389786 103254
rect 390022 103018 425786 103254
rect 426022 103018 461786 103254
rect 462022 103018 497786 103254
rect 498022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 591942 103254
rect 592178 103018 592360 103254
rect -8436 102934 592360 103018
rect -8436 102698 -8254 102934
rect -8018 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 317786 102934
rect 318022 102698 353786 102934
rect 354022 102698 389786 102934
rect 390022 102698 425786 102934
rect 426022 102698 461786 102934
rect 462022 102698 497786 102934
rect 498022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 591942 102934
rect 592178 102698 592360 102934
rect -8436 102676 592360 102698
rect -8436 102674 -7836 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 317604 102674 318204 102676
rect 353604 102674 354204 102676
rect 389604 102674 390204 102676
rect 425604 102674 426204 102676
rect 461604 102674 462204 102676
rect 497604 102674 498204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591760 102674 592360 102676
rect -6596 99676 -5996 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 589920 99676 590520 99678
rect -6596 99654 590520 99676
rect -6596 99418 -6414 99654
rect -6178 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590102 99654
rect 590338 99418 590520 99654
rect -6596 99334 590520 99418
rect -6596 99098 -6414 99334
rect -6178 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590102 99334
rect 590338 99098 590520 99334
rect -6596 99076 590520 99098
rect -6596 99074 -5996 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 589920 99074 590520 99076
rect -4756 96076 -4156 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588080 96076 588680 96078
rect -4756 96054 588680 96076
rect -4756 95818 -4574 96054
rect -4338 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588262 96054
rect 588498 95818 588680 96054
rect -4756 95734 588680 95818
rect -4756 95498 -4574 95734
rect -4338 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588262 95734
rect 588498 95498 588680 95734
rect -4756 95476 588680 95498
rect -4756 95474 -4156 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588080 95474 588680 95476
rect -2916 92476 -2316 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586240 92476 586840 92478
rect -2916 92454 586840 92476
rect -2916 92218 -2734 92454
rect -2498 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586422 92454
rect 586658 92218 586840 92454
rect -2916 92134 586840 92218
rect -2916 91898 -2734 92134
rect -2498 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586422 92134
rect 586658 91898 586840 92134
rect -2916 91876 586840 91898
rect -2916 91874 -2316 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586240 91874 586840 91876
rect -7516 85276 -6916 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590840 85276 591440 85278
rect -8436 85254 592360 85276
rect -8436 85018 -7334 85254
rect -7098 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591022 85254
rect 591258 85018 592360 85254
rect -8436 84934 592360 85018
rect -8436 84698 -7334 84934
rect -7098 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591022 84934
rect 591258 84698 592360 84934
rect -8436 84676 592360 84698
rect -7516 84674 -6916 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590840 84674 591440 84676
rect -5676 81676 -5076 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589000 81676 589600 81678
rect -6596 81654 590520 81676
rect -6596 81418 -5494 81654
rect -5258 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589182 81654
rect 589418 81418 590520 81654
rect -6596 81334 590520 81418
rect -6596 81098 -5494 81334
rect -5258 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589182 81334
rect 589418 81098 590520 81334
rect -6596 81076 590520 81098
rect -5676 81074 -5076 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589000 81074 589600 81076
rect -3836 78076 -3236 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587160 78076 587760 78078
rect -4756 78054 588680 78076
rect -4756 77818 -3654 78054
rect -3418 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587342 78054
rect 587578 77818 588680 78054
rect -4756 77734 588680 77818
rect -4756 77498 -3654 77734
rect -3418 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587342 77734
rect 587578 77498 588680 77734
rect -4756 77476 588680 77498
rect -3836 77474 -3236 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587160 77474 587760 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2916 74454 586840 74476
rect -2916 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586840 74454
rect -2916 74134 586840 74218
rect -2916 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586840 74134
rect -2916 73876 586840 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8436 67276 -7836 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591760 67276 592360 67278
rect -8436 67254 592360 67276
rect -8436 67018 -8254 67254
rect -8018 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 591942 67254
rect 592178 67018 592360 67254
rect -8436 66934 592360 67018
rect -8436 66698 -8254 66934
rect -8018 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 591942 66934
rect 592178 66698 592360 66934
rect -8436 66676 592360 66698
rect -8436 66674 -7836 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591760 66674 592360 66676
rect -6596 63676 -5996 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 589920 63676 590520 63678
rect -6596 63654 590520 63676
rect -6596 63418 -6414 63654
rect -6178 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590102 63654
rect 590338 63418 590520 63654
rect -6596 63334 590520 63418
rect -6596 63098 -6414 63334
rect -6178 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590102 63334
rect 590338 63098 590520 63334
rect -6596 63076 590520 63098
rect -6596 63074 -5996 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 589920 63074 590520 63076
rect -4756 60076 -4156 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588080 60076 588680 60078
rect -4756 60054 588680 60076
rect -4756 59818 -4574 60054
rect -4338 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588262 60054
rect 588498 59818 588680 60054
rect -4756 59734 588680 59818
rect -4756 59498 -4574 59734
rect -4338 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588262 59734
rect 588498 59498 588680 59734
rect -4756 59476 588680 59498
rect -4756 59474 -4156 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588080 59474 588680 59476
rect -2916 56476 -2316 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586240 56476 586840 56478
rect -2916 56454 586840 56476
rect -2916 56218 -2734 56454
rect -2498 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586422 56454
rect 586658 56218 586840 56454
rect -2916 56134 586840 56218
rect -2916 55898 -2734 56134
rect -2498 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586422 56134
rect 586658 55898 586840 56134
rect -2916 55876 586840 55898
rect -2916 55874 -2316 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586240 55874 586840 55876
rect -7516 49276 -6916 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590840 49276 591440 49278
rect -8436 49254 592360 49276
rect -8436 49018 -7334 49254
rect -7098 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591022 49254
rect 591258 49018 592360 49254
rect -8436 48934 592360 49018
rect -8436 48698 -7334 48934
rect -7098 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591022 48934
rect 591258 48698 592360 48934
rect -8436 48676 592360 48698
rect -7516 48674 -6916 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590840 48674 591440 48676
rect -5676 45676 -5076 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589000 45676 589600 45678
rect -6596 45654 590520 45676
rect -6596 45418 -5494 45654
rect -5258 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589182 45654
rect 589418 45418 590520 45654
rect -6596 45334 590520 45418
rect -6596 45098 -5494 45334
rect -5258 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589182 45334
rect 589418 45098 590520 45334
rect -6596 45076 590520 45098
rect -5676 45074 -5076 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589000 45074 589600 45076
rect -3836 42076 -3236 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587160 42076 587760 42078
rect -4756 42054 588680 42076
rect -4756 41818 -3654 42054
rect -3418 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587342 42054
rect 587578 41818 588680 42054
rect -4756 41734 588680 41818
rect -4756 41498 -3654 41734
rect -3418 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587342 41734
rect 587578 41498 588680 41734
rect -4756 41476 588680 41498
rect -3836 41474 -3236 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587160 41474 587760 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2916 38454 586840 38476
rect -2916 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586840 38454
rect -2916 38134 586840 38218
rect -2916 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586840 38134
rect -2916 37876 586840 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8436 31276 -7836 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591760 31276 592360 31278
rect -8436 31254 592360 31276
rect -8436 31018 -8254 31254
rect -8018 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 591942 31254
rect 592178 31018 592360 31254
rect -8436 30934 592360 31018
rect -8436 30698 -8254 30934
rect -8018 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 591942 30934
rect 592178 30698 592360 30934
rect -8436 30676 592360 30698
rect -8436 30674 -7836 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591760 30674 592360 30676
rect -6596 27676 -5996 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 589920 27676 590520 27678
rect -6596 27654 590520 27676
rect -6596 27418 -6414 27654
rect -6178 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590102 27654
rect 590338 27418 590520 27654
rect -6596 27334 590520 27418
rect -6596 27098 -6414 27334
rect -6178 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590102 27334
rect 590338 27098 590520 27334
rect -6596 27076 590520 27098
rect -6596 27074 -5996 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 589920 27074 590520 27076
rect -4756 24076 -4156 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588080 24076 588680 24078
rect -4756 24054 588680 24076
rect -4756 23818 -4574 24054
rect -4338 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588262 24054
rect 588498 23818 588680 24054
rect -4756 23734 588680 23818
rect -4756 23498 -4574 23734
rect -4338 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588262 23734
rect 588498 23498 588680 23734
rect -4756 23476 588680 23498
rect -4756 23474 -4156 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588080 23474 588680 23476
rect -2916 20476 -2316 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586240 20476 586840 20478
rect -2916 20454 586840 20476
rect -2916 20218 -2734 20454
rect -2498 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586422 20454
rect 586658 20218 586840 20454
rect -2916 20134 586840 20218
rect -2916 19898 -2734 20134
rect -2498 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586422 20134
rect 586658 19898 586840 20134
rect -2916 19876 586840 19898
rect -2916 19874 -2316 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586240 19874 586840 19876
rect -7516 13276 -6916 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590840 13276 591440 13278
rect -8436 13254 592360 13276
rect -8436 13018 -7334 13254
rect -7098 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591022 13254
rect 591258 13018 592360 13254
rect -8436 12934 592360 13018
rect -8436 12698 -7334 12934
rect -7098 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591022 12934
rect 591258 12698 592360 12934
rect -8436 12676 592360 12698
rect -7516 12674 -6916 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590840 12674 591440 12676
rect -5676 9676 -5076 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589000 9676 589600 9678
rect -6596 9654 590520 9676
rect -6596 9418 -5494 9654
rect -5258 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589182 9654
rect 589418 9418 590520 9654
rect -6596 9334 590520 9418
rect -6596 9098 -5494 9334
rect -5258 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589182 9334
rect 589418 9098 590520 9334
rect -6596 9076 590520 9098
rect -5676 9074 -5076 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589000 9074 589600 9076
rect -3836 6076 -3236 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587160 6076 587760 6078
rect -4756 6054 588680 6076
rect -4756 5818 -3654 6054
rect -3418 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587342 6054
rect 587578 5818 588680 6054
rect -4756 5734 588680 5818
rect -4756 5498 -3654 5734
rect -3418 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587342 5734
rect 587578 5498 588680 5734
rect -4756 5476 588680 5498
rect -3836 5474 -3236 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587160 5474 587760 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2916 2454 586840 2476
rect -2916 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586840 2454
rect -2916 2134 586840 2218
rect -2916 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586840 2134
rect -2916 1876 586840 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2916 -1244 -2316 -1242
rect 18804 -1244 19404 -1242
rect 54804 -1244 55404 -1242
rect 90804 -1244 91404 -1242
rect 126804 -1244 127404 -1242
rect 162804 -1244 163404 -1242
rect 198804 -1244 199404 -1242
rect 234804 -1244 235404 -1242
rect 270804 -1244 271404 -1242
rect 306804 -1244 307404 -1242
rect 342804 -1244 343404 -1242
rect 378804 -1244 379404 -1242
rect 414804 -1244 415404 -1242
rect 450804 -1244 451404 -1242
rect 486804 -1244 487404 -1242
rect 522804 -1244 523404 -1242
rect 558804 -1244 559404 -1242
rect 586240 -1244 586840 -1242
rect -2916 -1266 586840 -1244
rect -2916 -1502 -2734 -1266
rect -2498 -1502 18986 -1266
rect 19222 -1502 54986 -1266
rect 55222 -1502 90986 -1266
rect 91222 -1502 126986 -1266
rect 127222 -1502 162986 -1266
rect 163222 -1502 198986 -1266
rect 199222 -1502 234986 -1266
rect 235222 -1502 270986 -1266
rect 271222 -1502 306986 -1266
rect 307222 -1502 342986 -1266
rect 343222 -1502 378986 -1266
rect 379222 -1502 414986 -1266
rect 415222 -1502 450986 -1266
rect 451222 -1502 486986 -1266
rect 487222 -1502 522986 -1266
rect 523222 -1502 558986 -1266
rect 559222 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect -2916 -1586 586840 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 18986 -1586
rect 19222 -1822 54986 -1586
rect 55222 -1822 90986 -1586
rect 91222 -1822 126986 -1586
rect 127222 -1822 162986 -1586
rect 163222 -1822 198986 -1586
rect 199222 -1822 234986 -1586
rect 235222 -1822 270986 -1586
rect 271222 -1822 306986 -1586
rect 307222 -1822 342986 -1586
rect 343222 -1822 378986 -1586
rect 379222 -1822 414986 -1586
rect 415222 -1822 450986 -1586
rect 451222 -1822 486986 -1586
rect 487222 -1822 522986 -1586
rect 523222 -1822 558986 -1586
rect 559222 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect -2916 -1844 586840 -1822
rect -2916 -1846 -2316 -1844
rect 18804 -1846 19404 -1844
rect 54804 -1846 55404 -1844
rect 90804 -1846 91404 -1844
rect 126804 -1846 127404 -1844
rect 162804 -1846 163404 -1844
rect 198804 -1846 199404 -1844
rect 234804 -1846 235404 -1844
rect 270804 -1846 271404 -1844
rect 306804 -1846 307404 -1844
rect 342804 -1846 343404 -1844
rect 378804 -1846 379404 -1844
rect 414804 -1846 415404 -1844
rect 450804 -1846 451404 -1844
rect 486804 -1846 487404 -1844
rect 522804 -1846 523404 -1844
rect 558804 -1846 559404 -1844
rect 586240 -1846 586840 -1844
rect -3836 -2164 -3236 -2162
rect 4404 -2164 5004 -2162
rect 40404 -2164 41004 -2162
rect 76404 -2164 77004 -2162
rect 112404 -2164 113004 -2162
rect 148404 -2164 149004 -2162
rect 184404 -2164 185004 -2162
rect 220404 -2164 221004 -2162
rect 256404 -2164 257004 -2162
rect 292404 -2164 293004 -2162
rect 328404 -2164 329004 -2162
rect 364404 -2164 365004 -2162
rect 400404 -2164 401004 -2162
rect 436404 -2164 437004 -2162
rect 472404 -2164 473004 -2162
rect 508404 -2164 509004 -2162
rect 544404 -2164 545004 -2162
rect 580404 -2164 581004 -2162
rect 587160 -2164 587760 -2162
rect -3836 -2186 587760 -2164
rect -3836 -2422 -3654 -2186
rect -3418 -2422 4586 -2186
rect 4822 -2422 40586 -2186
rect 40822 -2422 76586 -2186
rect 76822 -2422 112586 -2186
rect 112822 -2422 148586 -2186
rect 148822 -2422 184586 -2186
rect 184822 -2422 220586 -2186
rect 220822 -2422 256586 -2186
rect 256822 -2422 292586 -2186
rect 292822 -2422 328586 -2186
rect 328822 -2422 364586 -2186
rect 364822 -2422 400586 -2186
rect 400822 -2422 436586 -2186
rect 436822 -2422 472586 -2186
rect 472822 -2422 508586 -2186
rect 508822 -2422 544586 -2186
rect 544822 -2422 580586 -2186
rect 580822 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect -3836 -2506 587760 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 4586 -2506
rect 4822 -2742 40586 -2506
rect 40822 -2742 76586 -2506
rect 76822 -2742 112586 -2506
rect 112822 -2742 148586 -2506
rect 148822 -2742 184586 -2506
rect 184822 -2742 220586 -2506
rect 220822 -2742 256586 -2506
rect 256822 -2742 292586 -2506
rect 292822 -2742 328586 -2506
rect 328822 -2742 364586 -2506
rect 364822 -2742 400586 -2506
rect 400822 -2742 436586 -2506
rect 436822 -2742 472586 -2506
rect 472822 -2742 508586 -2506
rect 508822 -2742 544586 -2506
rect 544822 -2742 580586 -2506
rect 580822 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect -3836 -2764 587760 -2742
rect -3836 -2766 -3236 -2764
rect 4404 -2766 5004 -2764
rect 40404 -2766 41004 -2764
rect 76404 -2766 77004 -2764
rect 112404 -2766 113004 -2764
rect 148404 -2766 149004 -2764
rect 184404 -2766 185004 -2764
rect 220404 -2766 221004 -2764
rect 256404 -2766 257004 -2764
rect 292404 -2766 293004 -2764
rect 328404 -2766 329004 -2764
rect 364404 -2766 365004 -2764
rect 400404 -2766 401004 -2764
rect 436404 -2766 437004 -2764
rect 472404 -2766 473004 -2764
rect 508404 -2766 509004 -2764
rect 544404 -2766 545004 -2764
rect 580404 -2766 581004 -2764
rect 587160 -2766 587760 -2764
rect -4756 -3084 -4156 -3082
rect 22404 -3084 23004 -3082
rect 58404 -3084 59004 -3082
rect 94404 -3084 95004 -3082
rect 130404 -3084 131004 -3082
rect 166404 -3084 167004 -3082
rect 202404 -3084 203004 -3082
rect 238404 -3084 239004 -3082
rect 274404 -3084 275004 -3082
rect 310404 -3084 311004 -3082
rect 346404 -3084 347004 -3082
rect 382404 -3084 383004 -3082
rect 418404 -3084 419004 -3082
rect 454404 -3084 455004 -3082
rect 490404 -3084 491004 -3082
rect 526404 -3084 527004 -3082
rect 562404 -3084 563004 -3082
rect 588080 -3084 588680 -3082
rect -4756 -3106 588680 -3084
rect -4756 -3342 -4574 -3106
rect -4338 -3342 22586 -3106
rect 22822 -3342 58586 -3106
rect 58822 -3342 94586 -3106
rect 94822 -3342 130586 -3106
rect 130822 -3342 166586 -3106
rect 166822 -3342 202586 -3106
rect 202822 -3342 238586 -3106
rect 238822 -3342 274586 -3106
rect 274822 -3342 310586 -3106
rect 310822 -3342 346586 -3106
rect 346822 -3342 382586 -3106
rect 382822 -3342 418586 -3106
rect 418822 -3342 454586 -3106
rect 454822 -3342 490586 -3106
rect 490822 -3342 526586 -3106
rect 526822 -3342 562586 -3106
rect 562822 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect -4756 -3426 588680 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 22586 -3426
rect 22822 -3662 58586 -3426
rect 58822 -3662 94586 -3426
rect 94822 -3662 130586 -3426
rect 130822 -3662 166586 -3426
rect 166822 -3662 202586 -3426
rect 202822 -3662 238586 -3426
rect 238822 -3662 274586 -3426
rect 274822 -3662 310586 -3426
rect 310822 -3662 346586 -3426
rect 346822 -3662 382586 -3426
rect 382822 -3662 418586 -3426
rect 418822 -3662 454586 -3426
rect 454822 -3662 490586 -3426
rect 490822 -3662 526586 -3426
rect 526822 -3662 562586 -3426
rect 562822 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect -4756 -3684 588680 -3662
rect -4756 -3686 -4156 -3684
rect 22404 -3686 23004 -3684
rect 58404 -3686 59004 -3684
rect 94404 -3686 95004 -3684
rect 130404 -3686 131004 -3684
rect 166404 -3686 167004 -3684
rect 202404 -3686 203004 -3684
rect 238404 -3686 239004 -3684
rect 274404 -3686 275004 -3684
rect 310404 -3686 311004 -3684
rect 346404 -3686 347004 -3684
rect 382404 -3686 383004 -3684
rect 418404 -3686 419004 -3684
rect 454404 -3686 455004 -3684
rect 490404 -3686 491004 -3684
rect 526404 -3686 527004 -3684
rect 562404 -3686 563004 -3684
rect 588080 -3686 588680 -3684
rect -5676 -4004 -5076 -4002
rect 8004 -4004 8604 -4002
rect 44004 -4004 44604 -4002
rect 80004 -4004 80604 -4002
rect 116004 -4004 116604 -4002
rect 152004 -4004 152604 -4002
rect 188004 -4004 188604 -4002
rect 224004 -4004 224604 -4002
rect 260004 -4004 260604 -4002
rect 296004 -4004 296604 -4002
rect 332004 -4004 332604 -4002
rect 368004 -4004 368604 -4002
rect 404004 -4004 404604 -4002
rect 440004 -4004 440604 -4002
rect 476004 -4004 476604 -4002
rect 512004 -4004 512604 -4002
rect 548004 -4004 548604 -4002
rect 589000 -4004 589600 -4002
rect -5676 -4026 589600 -4004
rect -5676 -4262 -5494 -4026
rect -5258 -4262 8186 -4026
rect 8422 -4262 44186 -4026
rect 44422 -4262 80186 -4026
rect 80422 -4262 116186 -4026
rect 116422 -4262 152186 -4026
rect 152422 -4262 188186 -4026
rect 188422 -4262 224186 -4026
rect 224422 -4262 260186 -4026
rect 260422 -4262 296186 -4026
rect 296422 -4262 332186 -4026
rect 332422 -4262 368186 -4026
rect 368422 -4262 404186 -4026
rect 404422 -4262 440186 -4026
rect 440422 -4262 476186 -4026
rect 476422 -4262 512186 -4026
rect 512422 -4262 548186 -4026
rect 548422 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect -5676 -4346 589600 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 8186 -4346
rect 8422 -4582 44186 -4346
rect 44422 -4582 80186 -4346
rect 80422 -4582 116186 -4346
rect 116422 -4582 152186 -4346
rect 152422 -4582 188186 -4346
rect 188422 -4582 224186 -4346
rect 224422 -4582 260186 -4346
rect 260422 -4582 296186 -4346
rect 296422 -4582 332186 -4346
rect 332422 -4582 368186 -4346
rect 368422 -4582 404186 -4346
rect 404422 -4582 440186 -4346
rect 440422 -4582 476186 -4346
rect 476422 -4582 512186 -4346
rect 512422 -4582 548186 -4346
rect 548422 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect -5676 -4604 589600 -4582
rect -5676 -4606 -5076 -4604
rect 8004 -4606 8604 -4604
rect 44004 -4606 44604 -4604
rect 80004 -4606 80604 -4604
rect 116004 -4606 116604 -4604
rect 152004 -4606 152604 -4604
rect 188004 -4606 188604 -4604
rect 224004 -4606 224604 -4604
rect 260004 -4606 260604 -4604
rect 296004 -4606 296604 -4604
rect 332004 -4606 332604 -4604
rect 368004 -4606 368604 -4604
rect 404004 -4606 404604 -4604
rect 440004 -4606 440604 -4604
rect 476004 -4606 476604 -4604
rect 512004 -4606 512604 -4604
rect 548004 -4606 548604 -4604
rect 589000 -4606 589600 -4604
rect -6596 -4924 -5996 -4922
rect 26004 -4924 26604 -4922
rect 62004 -4924 62604 -4922
rect 98004 -4924 98604 -4922
rect 134004 -4924 134604 -4922
rect 170004 -4924 170604 -4922
rect 206004 -4924 206604 -4922
rect 242004 -4924 242604 -4922
rect 278004 -4924 278604 -4922
rect 314004 -4924 314604 -4922
rect 350004 -4924 350604 -4922
rect 386004 -4924 386604 -4922
rect 422004 -4924 422604 -4922
rect 458004 -4924 458604 -4922
rect 494004 -4924 494604 -4922
rect 530004 -4924 530604 -4922
rect 566004 -4924 566604 -4922
rect 589920 -4924 590520 -4922
rect -6596 -4946 590520 -4924
rect -6596 -5182 -6414 -4946
rect -6178 -5182 26186 -4946
rect 26422 -5182 62186 -4946
rect 62422 -5182 98186 -4946
rect 98422 -5182 134186 -4946
rect 134422 -5182 170186 -4946
rect 170422 -5182 206186 -4946
rect 206422 -5182 242186 -4946
rect 242422 -5182 278186 -4946
rect 278422 -5182 314186 -4946
rect 314422 -5182 350186 -4946
rect 350422 -5182 386186 -4946
rect 386422 -5182 422186 -4946
rect 422422 -5182 458186 -4946
rect 458422 -5182 494186 -4946
rect 494422 -5182 530186 -4946
rect 530422 -5182 566186 -4946
rect 566422 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect -6596 -5266 590520 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 26186 -5266
rect 26422 -5502 62186 -5266
rect 62422 -5502 98186 -5266
rect 98422 -5502 134186 -5266
rect 134422 -5502 170186 -5266
rect 170422 -5502 206186 -5266
rect 206422 -5502 242186 -5266
rect 242422 -5502 278186 -5266
rect 278422 -5502 314186 -5266
rect 314422 -5502 350186 -5266
rect 350422 -5502 386186 -5266
rect 386422 -5502 422186 -5266
rect 422422 -5502 458186 -5266
rect 458422 -5502 494186 -5266
rect 494422 -5502 530186 -5266
rect 530422 -5502 566186 -5266
rect 566422 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect -6596 -5524 590520 -5502
rect -6596 -5526 -5996 -5524
rect 26004 -5526 26604 -5524
rect 62004 -5526 62604 -5524
rect 98004 -5526 98604 -5524
rect 134004 -5526 134604 -5524
rect 170004 -5526 170604 -5524
rect 206004 -5526 206604 -5524
rect 242004 -5526 242604 -5524
rect 278004 -5526 278604 -5524
rect 314004 -5526 314604 -5524
rect 350004 -5526 350604 -5524
rect 386004 -5526 386604 -5524
rect 422004 -5526 422604 -5524
rect 458004 -5526 458604 -5524
rect 494004 -5526 494604 -5524
rect 530004 -5526 530604 -5524
rect 566004 -5526 566604 -5524
rect 589920 -5526 590520 -5524
rect -7516 -5844 -6916 -5842
rect 11604 -5844 12204 -5842
rect 47604 -5844 48204 -5842
rect 83604 -5844 84204 -5842
rect 119604 -5844 120204 -5842
rect 155604 -5844 156204 -5842
rect 191604 -5844 192204 -5842
rect 227604 -5844 228204 -5842
rect 263604 -5844 264204 -5842
rect 299604 -5844 300204 -5842
rect 335604 -5844 336204 -5842
rect 371604 -5844 372204 -5842
rect 407604 -5844 408204 -5842
rect 443604 -5844 444204 -5842
rect 479604 -5844 480204 -5842
rect 515604 -5844 516204 -5842
rect 551604 -5844 552204 -5842
rect 590840 -5844 591440 -5842
rect -7516 -5866 591440 -5844
rect -7516 -6102 -7334 -5866
rect -7098 -6102 11786 -5866
rect 12022 -6102 47786 -5866
rect 48022 -6102 83786 -5866
rect 84022 -6102 119786 -5866
rect 120022 -6102 155786 -5866
rect 156022 -6102 191786 -5866
rect 192022 -6102 227786 -5866
rect 228022 -6102 263786 -5866
rect 264022 -6102 299786 -5866
rect 300022 -6102 335786 -5866
rect 336022 -6102 371786 -5866
rect 372022 -6102 407786 -5866
rect 408022 -6102 443786 -5866
rect 444022 -6102 479786 -5866
rect 480022 -6102 515786 -5866
rect 516022 -6102 551786 -5866
rect 552022 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect -7516 -6186 591440 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 11786 -6186
rect 12022 -6422 47786 -6186
rect 48022 -6422 83786 -6186
rect 84022 -6422 119786 -6186
rect 120022 -6422 155786 -6186
rect 156022 -6422 191786 -6186
rect 192022 -6422 227786 -6186
rect 228022 -6422 263786 -6186
rect 264022 -6422 299786 -6186
rect 300022 -6422 335786 -6186
rect 336022 -6422 371786 -6186
rect 372022 -6422 407786 -6186
rect 408022 -6422 443786 -6186
rect 444022 -6422 479786 -6186
rect 480022 -6422 515786 -6186
rect 516022 -6422 551786 -6186
rect 552022 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect -7516 -6444 591440 -6422
rect -7516 -6446 -6916 -6444
rect 11604 -6446 12204 -6444
rect 47604 -6446 48204 -6444
rect 83604 -6446 84204 -6444
rect 119604 -6446 120204 -6444
rect 155604 -6446 156204 -6444
rect 191604 -6446 192204 -6444
rect 227604 -6446 228204 -6444
rect 263604 -6446 264204 -6444
rect 299604 -6446 300204 -6444
rect 335604 -6446 336204 -6444
rect 371604 -6446 372204 -6444
rect 407604 -6446 408204 -6444
rect 443604 -6446 444204 -6444
rect 479604 -6446 480204 -6444
rect 515604 -6446 516204 -6444
rect 551604 -6446 552204 -6444
rect 590840 -6446 591440 -6444
rect -8436 -6764 -7836 -6762
rect 29604 -6764 30204 -6762
rect 65604 -6764 66204 -6762
rect 101604 -6764 102204 -6762
rect 137604 -6764 138204 -6762
rect 173604 -6764 174204 -6762
rect 209604 -6764 210204 -6762
rect 245604 -6764 246204 -6762
rect 281604 -6764 282204 -6762
rect 317604 -6764 318204 -6762
rect 353604 -6764 354204 -6762
rect 389604 -6764 390204 -6762
rect 425604 -6764 426204 -6762
rect 461604 -6764 462204 -6762
rect 497604 -6764 498204 -6762
rect 533604 -6764 534204 -6762
rect 569604 -6764 570204 -6762
rect 591760 -6764 592360 -6762
rect -8436 -6786 592360 -6764
rect -8436 -7022 -8254 -6786
rect -8018 -7022 29786 -6786
rect 30022 -7022 65786 -6786
rect 66022 -7022 101786 -6786
rect 102022 -7022 137786 -6786
rect 138022 -7022 173786 -6786
rect 174022 -7022 209786 -6786
rect 210022 -7022 245786 -6786
rect 246022 -7022 281786 -6786
rect 282022 -7022 317786 -6786
rect 318022 -7022 353786 -6786
rect 354022 -7022 389786 -6786
rect 390022 -7022 425786 -6786
rect 426022 -7022 461786 -6786
rect 462022 -7022 497786 -6786
rect 498022 -7022 533786 -6786
rect 534022 -7022 569786 -6786
rect 570022 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect -8436 -7106 592360 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 29786 -7106
rect 30022 -7342 65786 -7106
rect 66022 -7342 101786 -7106
rect 102022 -7342 137786 -7106
rect 138022 -7342 173786 -7106
rect 174022 -7342 209786 -7106
rect 210022 -7342 245786 -7106
rect 246022 -7342 281786 -7106
rect 282022 -7342 317786 -7106
rect 318022 -7342 353786 -7106
rect 354022 -7342 389786 -7106
rect 390022 -7342 425786 -7106
rect 426022 -7342 461786 -7106
rect 462022 -7342 497786 -7106
rect 498022 -7342 533786 -7106
rect 534022 -7342 569786 -7106
rect 570022 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect -8436 -7364 592360 -7342
rect -8436 -7366 -7836 -7364
rect 29604 -7366 30204 -7364
rect 65604 -7366 66204 -7364
rect 101604 -7366 102204 -7364
rect 137604 -7366 138204 -7364
rect 173604 -7366 174204 -7364
rect 209604 -7366 210204 -7364
rect 245604 -7366 246204 -7364
rect 281604 -7366 282204 -7364
rect 317604 -7366 318204 -7364
rect 353604 -7366 354204 -7364
rect 389604 -7366 390204 -7364
rect 425604 -7366 426204 -7364
rect 461604 -7366 462204 -7364
rect 497604 -7366 498204 -7364
rect 533604 -7366 534204 -7364
rect 569604 -7366 570204 -7364
rect 591760 -7366 592360 -7364
use user_proj_example  mprj
timestamp 1607074398
transform 1 0 230000 0 1 340000
box 0 0 119756 120000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 4 analog_io[0]
port 1 nsew
rlabel metal3 s 583520 474996 584960 475236 4 analog_io[10]
port 2 nsew
rlabel metal3 s 583520 521916 584960 522156 4 analog_io[11]
port 3 nsew
rlabel metal3 s 583520 568836 584960 569076 4 analog_io[12]
port 4 nsew
rlabel metal3 s 583520 615756 584960 615996 4 analog_io[13]
port 5 nsew
rlabel metal3 s 583520 662676 584960 662916 4 analog_io[14]
port 6 nsew
rlabel metal2 s 575818 703520 575930 704960 4 analog_io[15]
port 7 nsew
rlabel metal2 s 510958 703520 511070 704960 4 analog_io[16]
port 8 nsew
rlabel metal2 s 446098 703520 446210 704960 4 analog_io[17]
port 9 nsew
rlabel metal2 s 381146 703520 381258 704960 4 analog_io[18]
port 10 nsew
rlabel metal2 s 316286 703520 316398 704960 4 analog_io[19]
port 11 nsew
rlabel metal3 s 583520 52716 584960 52956 4 analog_io[1]
port 12 nsew
rlabel metal2 s 251426 703520 251538 704960 4 analog_io[20]
port 13 nsew
rlabel metal2 s 186474 703520 186586 704960 4 analog_io[21]
port 14 nsew
rlabel metal2 s 121614 703520 121726 704960 4 analog_io[22]
port 15 nsew
rlabel metal2 s 56754 703520 56866 704960 4 analog_io[23]
port 16 nsew
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 17 nsew
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 18 nsew
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 19 nsew
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 20 nsew
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 21 nsew
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 22 nsew
rlabel metal3 s 583520 99636 584960 99876 4 analog_io[2]
port 23 nsew
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 24 nsew
rlabel metal3 s 583520 146556 584960 146796 4 analog_io[3]
port 25 nsew
rlabel metal3 s 583520 193476 584960 193716 4 analog_io[4]
port 26 nsew
rlabel metal3 s 583520 240396 584960 240636 4 analog_io[5]
port 27 nsew
rlabel metal3 s 583520 287316 584960 287556 4 analog_io[6]
port 28 nsew
rlabel metal3 s 583520 334236 584960 334476 4 analog_io[7]
port 29 nsew
rlabel metal3 s 583520 381156 584960 381396 4 analog_io[8]
port 30 nsew
rlabel metal3 s 583520 428076 584960 428316 4 analog_io[9]
port 31 nsew
rlabel metal3 s 583520 17492 584960 17732 4 io_in[0]
port 32 nsew
rlabel metal3 s 583520 486692 584960 486932 4 io_in[10]
port 33 nsew
rlabel metal3 s 583520 533748 584960 533988 4 io_in[11]
port 34 nsew
rlabel metal3 s 583520 580668 584960 580908 4 io_in[12]
port 35 nsew
rlabel metal3 s 583520 627588 584960 627828 4 io_in[13]
port 36 nsew
rlabel metal3 s 583520 674508 584960 674748 4 io_in[14]
port 37 nsew
rlabel metal2 s 559626 703520 559738 704960 4 io_in[15]
port 38 nsew
rlabel metal2 s 494766 703520 494878 704960 4 io_in[16]
port 39 nsew
rlabel metal2 s 429814 703520 429926 704960 4 io_in[17]
port 40 nsew
rlabel metal2 s 364954 703520 365066 704960 4 io_in[18]
port 41 nsew
rlabel metal2 s 300094 703520 300206 704960 4 io_in[19]
port 42 nsew
rlabel metal3 s 583520 64412 584960 64652 4 io_in[1]
port 43 nsew
rlabel metal2 s 235142 703520 235254 704960 4 io_in[20]
port 44 nsew
rlabel metal2 s 170282 703520 170394 704960 4 io_in[21]
port 45 nsew
rlabel metal2 s 105422 703520 105534 704960 4 io_in[22]
port 46 nsew
rlabel metal2 s 40470 703520 40582 704960 4 io_in[23]
port 47 nsew
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 48 nsew
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 49 nsew
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 50 nsew
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 51 nsew
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 52 nsew
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 53 nsew
rlabel metal3 s 583520 111332 584960 111572 4 io_in[2]
port 54 nsew
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 55 nsew
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 56 nsew
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 57 nsew
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 58 nsew
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 59 nsew
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 60 nsew
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 61 nsew
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 62 nsew
rlabel metal3 s 583520 158252 584960 158492 4 io_in[3]
port 63 nsew
rlabel metal3 s 583520 205172 584960 205412 4 io_in[4]
port 64 nsew
rlabel metal3 s 583520 252092 584960 252332 4 io_in[5]
port 65 nsew
rlabel metal3 s 583520 299012 584960 299252 4 io_in[6]
port 66 nsew
rlabel metal3 s 583520 345932 584960 346172 4 io_in[7]
port 67 nsew
rlabel metal3 s 583520 392852 584960 393092 4 io_in[8]
port 68 nsew
rlabel metal3 s 583520 439772 584960 440012 4 io_in[9]
port 69 nsew
rlabel metal3 s 583520 40884 584960 41124 4 io_oeb[0]
port 70 nsew
rlabel metal3 s 583520 510220 584960 510460 4 io_oeb[10]
port 71 nsew
rlabel metal3 s 583520 557140 584960 557380 4 io_oeb[11]
port 72 nsew
rlabel metal3 s 583520 604060 584960 604300 4 io_oeb[12]
port 73 nsew
rlabel metal3 s 583520 650980 584960 651220 4 io_oeb[13]
port 74 nsew
rlabel metal3 s 583520 697900 584960 698140 4 io_oeb[14]
port 75 nsew
rlabel metal2 s 527150 703520 527262 704960 4 io_oeb[15]
port 76 nsew
rlabel metal2 s 462290 703520 462402 704960 4 io_oeb[16]
port 77 nsew
rlabel metal2 s 397430 703520 397542 704960 4 io_oeb[17]
port 78 nsew
rlabel metal2 s 332478 703520 332590 704960 4 io_oeb[18]
port 79 nsew
rlabel metal2 s 267618 703520 267730 704960 4 io_oeb[19]
port 80 nsew
rlabel metal3 s 583520 87804 584960 88044 4 io_oeb[1]
port 81 nsew
rlabel metal2 s 202758 703520 202870 704960 4 io_oeb[20]
port 82 nsew
rlabel metal2 s 137806 703520 137918 704960 4 io_oeb[21]
port 83 nsew
rlabel metal2 s 72946 703520 73058 704960 4 io_oeb[22]
port 84 nsew
rlabel metal2 s 8086 703520 8198 704960 4 io_oeb[23]
port 85 nsew
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 86 nsew
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 87 nsew
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 88 nsew
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 89 nsew
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 90 nsew
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 91 nsew
rlabel metal3 s 583520 134724 584960 134964 4 io_oeb[2]
port 92 nsew
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 93 nsew
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 94 nsew
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 95 nsew
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 96 nsew
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 97 nsew
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 98 nsew
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 99 nsew
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 100 nsew
rlabel metal3 s 583520 181780 584960 182020 4 io_oeb[3]
port 101 nsew
rlabel metal3 s 583520 228700 584960 228940 4 io_oeb[4]
port 102 nsew
rlabel metal3 s 583520 275620 584960 275860 4 io_oeb[5]
port 103 nsew
rlabel metal3 s 583520 322540 584960 322780 4 io_oeb[6]
port 104 nsew
rlabel metal3 s 583520 369460 584960 369700 4 io_oeb[7]
port 105 nsew
rlabel metal3 s 583520 416380 584960 416620 4 io_oeb[8]
port 106 nsew
rlabel metal3 s 583520 463300 584960 463540 4 io_oeb[9]
port 107 nsew
rlabel metal3 s 583520 29188 584960 29428 4 io_out[0]
port 108 nsew
rlabel metal3 s 583520 498524 584960 498764 4 io_out[10]
port 109 nsew
rlabel metal3 s 583520 545444 584960 545684 4 io_out[11]
port 110 nsew
rlabel metal3 s 583520 592364 584960 592604 4 io_out[12]
port 111 nsew
rlabel metal3 s 583520 639284 584960 639524 4 io_out[13]
port 112 nsew
rlabel metal3 s 583520 686204 584960 686444 4 io_out[14]
port 113 nsew
rlabel metal2 s 543434 703520 543546 704960 4 io_out[15]
port 114 nsew
rlabel metal2 s 478482 703520 478594 704960 4 io_out[16]
port 115 nsew
rlabel metal2 s 413622 703520 413734 704960 4 io_out[17]
port 116 nsew
rlabel metal2 s 348762 703520 348874 704960 4 io_out[18]
port 117 nsew
rlabel metal2 s 283810 703520 283922 704960 4 io_out[19]
port 118 nsew
rlabel metal3 s 583520 76108 584960 76348 4 io_out[1]
port 119 nsew
rlabel metal2 s 218950 703520 219062 704960 4 io_out[20]
port 120 nsew
rlabel metal2 s 154090 703520 154202 704960 4 io_out[21]
port 121 nsew
rlabel metal2 s 89138 703520 89250 704960 4 io_out[22]
port 122 nsew
rlabel metal2 s 24278 703520 24390 704960 4 io_out[23]
port 123 nsew
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 124 nsew
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 125 nsew
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 126 nsew
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 127 nsew
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 128 nsew
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 129 nsew
rlabel metal3 s 583520 123028 584960 123268 4 io_out[2]
port 130 nsew
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 131 nsew
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 132 nsew
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 133 nsew
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 134 nsew
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 135 nsew
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 136 nsew
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 137 nsew
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 138 nsew
rlabel metal3 s 583520 169948 584960 170188 4 io_out[3]
port 139 nsew
rlabel metal3 s 583520 216868 584960 217108 4 io_out[4]
port 140 nsew
rlabel metal3 s 583520 263788 584960 264028 4 io_out[5]
port 141 nsew
rlabel metal3 s 583520 310708 584960 310948 4 io_out[6]
port 142 nsew
rlabel metal3 s 583520 357764 584960 358004 4 io_out[7]
port 143 nsew
rlabel metal3 s 583520 404684 584960 404924 4 io_out[8]
port 144 nsew
rlabel metal3 s 583520 451604 584960 451844 4 io_out[9]
port 145 nsew
rlabel metal2 s 126582 -960 126694 480 4 la_data_in[0]
port 146 nsew
rlabel metal2 s 483450 -960 483562 480 4 la_data_in[100]
port 147 nsew
rlabel metal2 s 486946 -960 487058 480 4 la_data_in[101]
port 148 nsew
rlabel metal2 s 490534 -960 490646 480 4 la_data_in[102]
port 149 nsew
rlabel metal2 s 494122 -960 494234 480 4 la_data_in[103]
port 150 nsew
rlabel metal2 s 497710 -960 497822 480 4 la_data_in[104]
port 151 nsew
rlabel metal2 s 501206 -960 501318 480 4 la_data_in[105]
port 152 nsew
rlabel metal2 s 504794 -960 504906 480 4 la_data_in[106]
port 153 nsew
rlabel metal2 s 508382 -960 508494 480 4 la_data_in[107]
port 154 nsew
rlabel metal2 s 511970 -960 512082 480 4 la_data_in[108]
port 155 nsew
rlabel metal2 s 515558 -960 515670 480 4 la_data_in[109]
port 156 nsew
rlabel metal2 s 162278 -960 162390 480 4 la_data_in[10]
port 157 nsew
rlabel metal2 s 519054 -960 519166 480 4 la_data_in[110]
port 158 nsew
rlabel metal2 s 522642 -960 522754 480 4 la_data_in[111]
port 159 nsew
rlabel metal2 s 526230 -960 526342 480 4 la_data_in[112]
port 160 nsew
rlabel metal2 s 529818 -960 529930 480 4 la_data_in[113]
port 161 nsew
rlabel metal2 s 533406 -960 533518 480 4 la_data_in[114]
port 162 nsew
rlabel metal2 s 536902 -960 537014 480 4 la_data_in[115]
port 163 nsew
rlabel metal2 s 540490 -960 540602 480 4 la_data_in[116]
port 164 nsew
rlabel metal2 s 544078 -960 544190 480 4 la_data_in[117]
port 165 nsew
rlabel metal2 s 547666 -960 547778 480 4 la_data_in[118]
port 166 nsew
rlabel metal2 s 551162 -960 551274 480 4 la_data_in[119]
port 167 nsew
rlabel metal2 s 165866 -960 165978 480 4 la_data_in[11]
port 168 nsew
rlabel metal2 s 554750 -960 554862 480 4 la_data_in[120]
port 169 nsew
rlabel metal2 s 558338 -960 558450 480 4 la_data_in[121]
port 170 nsew
rlabel metal2 s 561926 -960 562038 480 4 la_data_in[122]
port 171 nsew
rlabel metal2 s 565514 -960 565626 480 4 la_data_in[123]
port 172 nsew
rlabel metal2 s 569010 -960 569122 480 4 la_data_in[124]
port 173 nsew
rlabel metal2 s 572598 -960 572710 480 4 la_data_in[125]
port 174 nsew
rlabel metal2 s 576186 -960 576298 480 4 la_data_in[126]
port 175 nsew
rlabel metal2 s 579774 -960 579886 480 4 la_data_in[127]
port 176 nsew
rlabel metal2 s 169362 -960 169474 480 4 la_data_in[12]
port 177 nsew
rlabel metal2 s 172950 -960 173062 480 4 la_data_in[13]
port 178 nsew
rlabel metal2 s 176538 -960 176650 480 4 la_data_in[14]
port 179 nsew
rlabel metal2 s 180126 -960 180238 480 4 la_data_in[15]
port 180 nsew
rlabel metal2 s 183714 -960 183826 480 4 la_data_in[16]
port 181 nsew
rlabel metal2 s 187210 -960 187322 480 4 la_data_in[17]
port 182 nsew
rlabel metal2 s 190798 -960 190910 480 4 la_data_in[18]
port 183 nsew
rlabel metal2 s 194386 -960 194498 480 4 la_data_in[19]
port 184 nsew
rlabel metal2 s 130170 -960 130282 480 4 la_data_in[1]
port 185 nsew
rlabel metal2 s 197974 -960 198086 480 4 la_data_in[20]
port 186 nsew
rlabel metal2 s 201470 -960 201582 480 4 la_data_in[21]
port 187 nsew
rlabel metal2 s 205058 -960 205170 480 4 la_data_in[22]
port 188 nsew
rlabel metal2 s 208646 -960 208758 480 4 la_data_in[23]
port 189 nsew
rlabel metal2 s 212234 -960 212346 480 4 la_data_in[24]
port 190 nsew
rlabel metal2 s 215822 -960 215934 480 4 la_data_in[25]
port 191 nsew
rlabel metal2 s 219318 -960 219430 480 4 la_data_in[26]
port 192 nsew
rlabel metal2 s 222906 -960 223018 480 4 la_data_in[27]
port 193 nsew
rlabel metal2 s 226494 -960 226606 480 4 la_data_in[28]
port 194 nsew
rlabel metal2 s 230082 -960 230194 480 4 la_data_in[29]
port 195 nsew
rlabel metal2 s 133758 -960 133870 480 4 la_data_in[2]
port 196 nsew
rlabel metal2 s 233670 -960 233782 480 4 la_data_in[30]
port 197 nsew
rlabel metal2 s 237166 -960 237278 480 4 la_data_in[31]
port 198 nsew
rlabel metal2 s 240754 -960 240866 480 4 la_data_in[32]
port 199 nsew
rlabel metal2 s 244342 -960 244454 480 4 la_data_in[33]
port 200 nsew
rlabel metal2 s 247930 -960 248042 480 4 la_data_in[34]
port 201 nsew
rlabel metal2 s 251426 -960 251538 480 4 la_data_in[35]
port 202 nsew
rlabel metal2 s 255014 -960 255126 480 4 la_data_in[36]
port 203 nsew
rlabel metal2 s 258602 -960 258714 480 4 la_data_in[37]
port 204 nsew
rlabel metal2 s 262190 -960 262302 480 4 la_data_in[38]
port 205 nsew
rlabel metal2 s 265778 -960 265890 480 4 la_data_in[39]
port 206 nsew
rlabel metal2 s 137254 -960 137366 480 4 la_data_in[3]
port 207 nsew
rlabel metal2 s 269274 -960 269386 480 4 la_data_in[40]
port 208 nsew
rlabel metal2 s 272862 -960 272974 480 4 la_data_in[41]
port 209 nsew
rlabel metal2 s 276450 -960 276562 480 4 la_data_in[42]
port 210 nsew
rlabel metal2 s 280038 -960 280150 480 4 la_data_in[43]
port 211 nsew
rlabel metal2 s 283626 -960 283738 480 4 la_data_in[44]
port 212 nsew
rlabel metal2 s 287122 -960 287234 480 4 la_data_in[45]
port 213 nsew
rlabel metal2 s 290710 -960 290822 480 4 la_data_in[46]
port 214 nsew
rlabel metal2 s 294298 -960 294410 480 4 la_data_in[47]
port 215 nsew
rlabel metal2 s 297886 -960 297998 480 4 la_data_in[48]
port 216 nsew
rlabel metal2 s 301382 -960 301494 480 4 la_data_in[49]
port 217 nsew
rlabel metal2 s 140842 -960 140954 480 4 la_data_in[4]
port 218 nsew
rlabel metal2 s 304970 -960 305082 480 4 la_data_in[50]
port 219 nsew
rlabel metal2 s 308558 -960 308670 480 4 la_data_in[51]
port 220 nsew
rlabel metal2 s 312146 -960 312258 480 4 la_data_in[52]
port 221 nsew
rlabel metal2 s 315734 -960 315846 480 4 la_data_in[53]
port 222 nsew
rlabel metal2 s 319230 -960 319342 480 4 la_data_in[54]
port 223 nsew
rlabel metal2 s 322818 -960 322930 480 4 la_data_in[55]
port 224 nsew
rlabel metal2 s 326406 -960 326518 480 4 la_data_in[56]
port 225 nsew
rlabel metal2 s 329994 -960 330106 480 4 la_data_in[57]
port 226 nsew
rlabel metal2 s 333582 -960 333694 480 4 la_data_in[58]
port 227 nsew
rlabel metal2 s 337078 -960 337190 480 4 la_data_in[59]
port 228 nsew
rlabel metal2 s 144430 -960 144542 480 4 la_data_in[5]
port 229 nsew
rlabel metal2 s 340666 -960 340778 480 4 la_data_in[60]
port 230 nsew
rlabel metal2 s 344254 -960 344366 480 4 la_data_in[61]
port 231 nsew
rlabel metal2 s 347842 -960 347954 480 4 la_data_in[62]
port 232 nsew
rlabel metal2 s 351338 -960 351450 480 4 la_data_in[63]
port 233 nsew
rlabel metal2 s 354926 -960 355038 480 4 la_data_in[64]
port 234 nsew
rlabel metal2 s 358514 -960 358626 480 4 la_data_in[65]
port 235 nsew
rlabel metal2 s 362102 -960 362214 480 4 la_data_in[66]
port 236 nsew
rlabel metal2 s 365690 -960 365802 480 4 la_data_in[67]
port 237 nsew
rlabel metal2 s 369186 -960 369298 480 4 la_data_in[68]
port 238 nsew
rlabel metal2 s 372774 -960 372886 480 4 la_data_in[69]
port 239 nsew
rlabel metal2 s 148018 -960 148130 480 4 la_data_in[6]
port 240 nsew
rlabel metal2 s 376362 -960 376474 480 4 la_data_in[70]
port 241 nsew
rlabel metal2 s 379950 -960 380062 480 4 la_data_in[71]
port 242 nsew
rlabel metal2 s 383538 -960 383650 480 4 la_data_in[72]
port 243 nsew
rlabel metal2 s 387034 -960 387146 480 4 la_data_in[73]
port 244 nsew
rlabel metal2 s 390622 -960 390734 480 4 la_data_in[74]
port 245 nsew
rlabel metal2 s 394210 -960 394322 480 4 la_data_in[75]
port 246 nsew
rlabel metal2 s 397798 -960 397910 480 4 la_data_in[76]
port 247 nsew
rlabel metal2 s 401294 -960 401406 480 4 la_data_in[77]
port 248 nsew
rlabel metal2 s 404882 -960 404994 480 4 la_data_in[78]
port 249 nsew
rlabel metal2 s 408470 -960 408582 480 4 la_data_in[79]
port 250 nsew
rlabel metal2 s 151514 -960 151626 480 4 la_data_in[7]
port 251 nsew
rlabel metal2 s 412058 -960 412170 480 4 la_data_in[80]
port 252 nsew
rlabel metal2 s 415646 -960 415758 480 4 la_data_in[81]
port 253 nsew
rlabel metal2 s 419142 -960 419254 480 4 la_data_in[82]
port 254 nsew
rlabel metal2 s 422730 -960 422842 480 4 la_data_in[83]
port 255 nsew
rlabel metal2 s 426318 -960 426430 480 4 la_data_in[84]
port 256 nsew
rlabel metal2 s 429906 -960 430018 480 4 la_data_in[85]
port 257 nsew
rlabel metal2 s 433494 -960 433606 480 4 la_data_in[86]
port 258 nsew
rlabel metal2 s 436990 -960 437102 480 4 la_data_in[87]
port 259 nsew
rlabel metal2 s 440578 -960 440690 480 4 la_data_in[88]
port 260 nsew
rlabel metal2 s 444166 -960 444278 480 4 la_data_in[89]
port 261 nsew
rlabel metal2 s 155102 -960 155214 480 4 la_data_in[8]
port 262 nsew
rlabel metal2 s 447754 -960 447866 480 4 la_data_in[90]
port 263 nsew
rlabel metal2 s 451250 -960 451362 480 4 la_data_in[91]
port 264 nsew
rlabel metal2 s 454838 -960 454950 480 4 la_data_in[92]
port 265 nsew
rlabel metal2 s 458426 -960 458538 480 4 la_data_in[93]
port 266 nsew
rlabel metal2 s 462014 -960 462126 480 4 la_data_in[94]
port 267 nsew
rlabel metal2 s 465602 -960 465714 480 4 la_data_in[95]
port 268 nsew
rlabel metal2 s 469098 -960 469210 480 4 la_data_in[96]
port 269 nsew
rlabel metal2 s 472686 -960 472798 480 4 la_data_in[97]
port 270 nsew
rlabel metal2 s 476274 -960 476386 480 4 la_data_in[98]
port 271 nsew
rlabel metal2 s 479862 -960 479974 480 4 la_data_in[99]
port 272 nsew
rlabel metal2 s 158690 -960 158802 480 4 la_data_in[9]
port 273 nsew
rlabel metal2 s 127778 -960 127890 480 4 la_data_out[0]
port 274 nsew
rlabel metal2 s 484554 -960 484666 480 4 la_data_out[100]
port 275 nsew
rlabel metal2 s 488142 -960 488254 480 4 la_data_out[101]
port 276 nsew
rlabel metal2 s 491730 -960 491842 480 4 la_data_out[102]
port 277 nsew
rlabel metal2 s 495318 -960 495430 480 4 la_data_out[103]
port 278 nsew
rlabel metal2 s 498906 -960 499018 480 4 la_data_out[104]
port 279 nsew
rlabel metal2 s 502402 -960 502514 480 4 la_data_out[105]
port 280 nsew
rlabel metal2 s 505990 -960 506102 480 4 la_data_out[106]
port 281 nsew
rlabel metal2 s 509578 -960 509690 480 4 la_data_out[107]
port 282 nsew
rlabel metal2 s 513166 -960 513278 480 4 la_data_out[108]
port 283 nsew
rlabel metal2 s 516754 -960 516866 480 4 la_data_out[109]
port 284 nsew
rlabel metal2 s 163474 -960 163586 480 4 la_data_out[10]
port 285 nsew
rlabel metal2 s 520250 -960 520362 480 4 la_data_out[110]
port 286 nsew
rlabel metal2 s 523838 -960 523950 480 4 la_data_out[111]
port 287 nsew
rlabel metal2 s 527426 -960 527538 480 4 la_data_out[112]
port 288 nsew
rlabel metal2 s 531014 -960 531126 480 4 la_data_out[113]
port 289 nsew
rlabel metal2 s 534510 -960 534622 480 4 la_data_out[114]
port 290 nsew
rlabel metal2 s 538098 -960 538210 480 4 la_data_out[115]
port 291 nsew
rlabel metal2 s 541686 -960 541798 480 4 la_data_out[116]
port 292 nsew
rlabel metal2 s 545274 -960 545386 480 4 la_data_out[117]
port 293 nsew
rlabel metal2 s 548862 -960 548974 480 4 la_data_out[118]
port 294 nsew
rlabel metal2 s 552358 -960 552470 480 4 la_data_out[119]
port 295 nsew
rlabel metal2 s 167062 -960 167174 480 4 la_data_out[11]
port 296 nsew
rlabel metal2 s 555946 -960 556058 480 4 la_data_out[120]
port 297 nsew
rlabel metal2 s 559534 -960 559646 480 4 la_data_out[121]
port 298 nsew
rlabel metal2 s 563122 -960 563234 480 4 la_data_out[122]
port 299 nsew
rlabel metal2 s 566710 -960 566822 480 4 la_data_out[123]
port 300 nsew
rlabel metal2 s 570206 -960 570318 480 4 la_data_out[124]
port 301 nsew
rlabel metal2 s 573794 -960 573906 480 4 la_data_out[125]
port 302 nsew
rlabel metal2 s 577382 -960 577494 480 4 la_data_out[126]
port 303 nsew
rlabel metal2 s 580970 -960 581082 480 4 la_data_out[127]
port 304 nsew
rlabel metal2 s 170558 -960 170670 480 4 la_data_out[12]
port 305 nsew
rlabel metal2 s 174146 -960 174258 480 4 la_data_out[13]
port 306 nsew
rlabel metal2 s 177734 -960 177846 480 4 la_data_out[14]
port 307 nsew
rlabel metal2 s 181322 -960 181434 480 4 la_data_out[15]
port 308 nsew
rlabel metal2 s 184818 -960 184930 480 4 la_data_out[16]
port 309 nsew
rlabel metal2 s 188406 -960 188518 480 4 la_data_out[17]
port 310 nsew
rlabel metal2 s 191994 -960 192106 480 4 la_data_out[18]
port 311 nsew
rlabel metal2 s 195582 -960 195694 480 4 la_data_out[19]
port 312 nsew
rlabel metal2 s 131366 -960 131478 480 4 la_data_out[1]
port 313 nsew
rlabel metal2 s 199170 -960 199282 480 4 la_data_out[20]
port 314 nsew
rlabel metal2 s 202666 -960 202778 480 4 la_data_out[21]
port 315 nsew
rlabel metal2 s 206254 -960 206366 480 4 la_data_out[22]
port 316 nsew
rlabel metal2 s 209842 -960 209954 480 4 la_data_out[23]
port 317 nsew
rlabel metal2 s 213430 -960 213542 480 4 la_data_out[24]
port 318 nsew
rlabel metal2 s 217018 -960 217130 480 4 la_data_out[25]
port 319 nsew
rlabel metal2 s 220514 -960 220626 480 4 la_data_out[26]
port 320 nsew
rlabel metal2 s 224102 -960 224214 480 4 la_data_out[27]
port 321 nsew
rlabel metal2 s 227690 -960 227802 480 4 la_data_out[28]
port 322 nsew
rlabel metal2 s 231278 -960 231390 480 4 la_data_out[29]
port 323 nsew
rlabel metal2 s 134862 -960 134974 480 4 la_data_out[2]
port 324 nsew
rlabel metal2 s 234774 -960 234886 480 4 la_data_out[30]
port 325 nsew
rlabel metal2 s 238362 -960 238474 480 4 la_data_out[31]
port 326 nsew
rlabel metal2 s 241950 -960 242062 480 4 la_data_out[32]
port 327 nsew
rlabel metal2 s 245538 -960 245650 480 4 la_data_out[33]
port 328 nsew
rlabel metal2 s 249126 -960 249238 480 4 la_data_out[34]
port 329 nsew
rlabel metal2 s 252622 -960 252734 480 4 la_data_out[35]
port 330 nsew
rlabel metal2 s 256210 -960 256322 480 4 la_data_out[36]
port 331 nsew
rlabel metal2 s 259798 -960 259910 480 4 la_data_out[37]
port 332 nsew
rlabel metal2 s 263386 -960 263498 480 4 la_data_out[38]
port 333 nsew
rlabel metal2 s 266974 -960 267086 480 4 la_data_out[39]
port 334 nsew
rlabel metal2 s 138450 -960 138562 480 4 la_data_out[3]
port 335 nsew
rlabel metal2 s 270470 -960 270582 480 4 la_data_out[40]
port 336 nsew
rlabel metal2 s 274058 -960 274170 480 4 la_data_out[41]
port 337 nsew
rlabel metal2 s 277646 -960 277758 480 4 la_data_out[42]
port 338 nsew
rlabel metal2 s 281234 -960 281346 480 4 la_data_out[43]
port 339 nsew
rlabel metal2 s 284730 -960 284842 480 4 la_data_out[44]
port 340 nsew
rlabel metal2 s 288318 -960 288430 480 4 la_data_out[45]
port 341 nsew
rlabel metal2 s 291906 -960 292018 480 4 la_data_out[46]
port 342 nsew
rlabel metal2 s 295494 -960 295606 480 4 la_data_out[47]
port 343 nsew
rlabel metal2 s 299082 -960 299194 480 4 la_data_out[48]
port 344 nsew
rlabel metal2 s 302578 -960 302690 480 4 la_data_out[49]
port 345 nsew
rlabel metal2 s 142038 -960 142150 480 4 la_data_out[4]
port 346 nsew
rlabel metal2 s 306166 -960 306278 480 4 la_data_out[50]
port 347 nsew
rlabel metal2 s 309754 -960 309866 480 4 la_data_out[51]
port 348 nsew
rlabel metal2 s 313342 -960 313454 480 4 la_data_out[52]
port 349 nsew
rlabel metal2 s 316930 -960 317042 480 4 la_data_out[53]
port 350 nsew
rlabel metal2 s 320426 -960 320538 480 4 la_data_out[54]
port 351 nsew
rlabel metal2 s 324014 -960 324126 480 4 la_data_out[55]
port 352 nsew
rlabel metal2 s 327602 -960 327714 480 4 la_data_out[56]
port 353 nsew
rlabel metal2 s 331190 -960 331302 480 4 la_data_out[57]
port 354 nsew
rlabel metal2 s 334686 -960 334798 480 4 la_data_out[58]
port 355 nsew
rlabel metal2 s 338274 -960 338386 480 4 la_data_out[59]
port 356 nsew
rlabel metal2 s 145626 -960 145738 480 4 la_data_out[5]
port 357 nsew
rlabel metal2 s 341862 -960 341974 480 4 la_data_out[60]
port 358 nsew
rlabel metal2 s 345450 -960 345562 480 4 la_data_out[61]
port 359 nsew
rlabel metal2 s 349038 -960 349150 480 4 la_data_out[62]
port 360 nsew
rlabel metal2 s 352534 -960 352646 480 4 la_data_out[63]
port 361 nsew
rlabel metal2 s 356122 -960 356234 480 4 la_data_out[64]
port 362 nsew
rlabel metal2 s 359710 -960 359822 480 4 la_data_out[65]
port 363 nsew
rlabel metal2 s 363298 -960 363410 480 4 la_data_out[66]
port 364 nsew
rlabel metal2 s 366886 -960 366998 480 4 la_data_out[67]
port 365 nsew
rlabel metal2 s 370382 -960 370494 480 4 la_data_out[68]
port 366 nsew
rlabel metal2 s 373970 -960 374082 480 4 la_data_out[69]
port 367 nsew
rlabel metal2 s 149214 -960 149326 480 4 la_data_out[6]
port 368 nsew
rlabel metal2 s 377558 -960 377670 480 4 la_data_out[70]
port 369 nsew
rlabel metal2 s 381146 -960 381258 480 4 la_data_out[71]
port 370 nsew
rlabel metal2 s 384642 -960 384754 480 4 la_data_out[72]
port 371 nsew
rlabel metal2 s 388230 -960 388342 480 4 la_data_out[73]
port 372 nsew
rlabel metal2 s 391818 -960 391930 480 4 la_data_out[74]
port 373 nsew
rlabel metal2 s 395406 -960 395518 480 4 la_data_out[75]
port 374 nsew
rlabel metal2 s 398994 -960 399106 480 4 la_data_out[76]
port 375 nsew
rlabel metal2 s 402490 -960 402602 480 4 la_data_out[77]
port 376 nsew
rlabel metal2 s 406078 -960 406190 480 4 la_data_out[78]
port 377 nsew
rlabel metal2 s 409666 -960 409778 480 4 la_data_out[79]
port 378 nsew
rlabel metal2 s 152710 -960 152822 480 4 la_data_out[7]
port 379 nsew
rlabel metal2 s 413254 -960 413366 480 4 la_data_out[80]
port 380 nsew
rlabel metal2 s 416842 -960 416954 480 4 la_data_out[81]
port 381 nsew
rlabel metal2 s 420338 -960 420450 480 4 la_data_out[82]
port 382 nsew
rlabel metal2 s 423926 -960 424038 480 4 la_data_out[83]
port 383 nsew
rlabel metal2 s 427514 -960 427626 480 4 la_data_out[84]
port 384 nsew
rlabel metal2 s 431102 -960 431214 480 4 la_data_out[85]
port 385 nsew
rlabel metal2 s 434598 -960 434710 480 4 la_data_out[86]
port 386 nsew
rlabel metal2 s 438186 -960 438298 480 4 la_data_out[87]
port 387 nsew
rlabel metal2 s 441774 -960 441886 480 4 la_data_out[88]
port 388 nsew
rlabel metal2 s 445362 -960 445474 480 4 la_data_out[89]
port 389 nsew
rlabel metal2 s 156298 -960 156410 480 4 la_data_out[8]
port 390 nsew
rlabel metal2 s 448950 -960 449062 480 4 la_data_out[90]
port 391 nsew
rlabel metal2 s 452446 -960 452558 480 4 la_data_out[91]
port 392 nsew
rlabel metal2 s 456034 -960 456146 480 4 la_data_out[92]
port 393 nsew
rlabel metal2 s 459622 -960 459734 480 4 la_data_out[93]
port 394 nsew
rlabel metal2 s 463210 -960 463322 480 4 la_data_out[94]
port 395 nsew
rlabel metal2 s 466798 -960 466910 480 4 la_data_out[95]
port 396 nsew
rlabel metal2 s 470294 -960 470406 480 4 la_data_out[96]
port 397 nsew
rlabel metal2 s 473882 -960 473994 480 4 la_data_out[97]
port 398 nsew
rlabel metal2 s 477470 -960 477582 480 4 la_data_out[98]
port 399 nsew
rlabel metal2 s 481058 -960 481170 480 4 la_data_out[99]
port 400 nsew
rlabel metal2 s 159886 -960 159998 480 4 la_data_out[9]
port 401 nsew
rlabel metal2 s 128974 -960 129086 480 4 la_oen[0]
port 402 nsew
rlabel metal2 s 485750 -960 485862 480 4 la_oen[100]
port 403 nsew
rlabel metal2 s 489338 -960 489450 480 4 la_oen[101]
port 404 nsew
rlabel metal2 s 492926 -960 493038 480 4 la_oen[102]
port 405 nsew
rlabel metal2 s 496514 -960 496626 480 4 la_oen[103]
port 406 nsew
rlabel metal2 s 500102 -960 500214 480 4 la_oen[104]
port 407 nsew
rlabel metal2 s 503598 -960 503710 480 4 la_oen[105]
port 408 nsew
rlabel metal2 s 507186 -960 507298 480 4 la_oen[106]
port 409 nsew
rlabel metal2 s 510774 -960 510886 480 4 la_oen[107]
port 410 nsew
rlabel metal2 s 514362 -960 514474 480 4 la_oen[108]
port 411 nsew
rlabel metal2 s 517858 -960 517970 480 4 la_oen[109]
port 412 nsew
rlabel metal2 s 164670 -960 164782 480 4 la_oen[10]
port 413 nsew
rlabel metal2 s 521446 -960 521558 480 4 la_oen[110]
port 414 nsew
rlabel metal2 s 525034 -960 525146 480 4 la_oen[111]
port 415 nsew
rlabel metal2 s 528622 -960 528734 480 4 la_oen[112]
port 416 nsew
rlabel metal2 s 532210 -960 532322 480 4 la_oen[113]
port 417 nsew
rlabel metal2 s 535706 -960 535818 480 4 la_oen[114]
port 418 nsew
rlabel metal2 s 539294 -960 539406 480 4 la_oen[115]
port 419 nsew
rlabel metal2 s 542882 -960 542994 480 4 la_oen[116]
port 420 nsew
rlabel metal2 s 546470 -960 546582 480 4 la_oen[117]
port 421 nsew
rlabel metal2 s 550058 -960 550170 480 4 la_oen[118]
port 422 nsew
rlabel metal2 s 553554 -960 553666 480 4 la_oen[119]
port 423 nsew
rlabel metal2 s 168166 -960 168278 480 4 la_oen[11]
port 424 nsew
rlabel metal2 s 557142 -960 557254 480 4 la_oen[120]
port 425 nsew
rlabel metal2 s 560730 -960 560842 480 4 la_oen[121]
port 426 nsew
rlabel metal2 s 564318 -960 564430 480 4 la_oen[122]
port 427 nsew
rlabel metal2 s 567814 -960 567926 480 4 la_oen[123]
port 428 nsew
rlabel metal2 s 571402 -960 571514 480 4 la_oen[124]
port 429 nsew
rlabel metal2 s 574990 -960 575102 480 4 la_oen[125]
port 430 nsew
rlabel metal2 s 578578 -960 578690 480 4 la_oen[126]
port 431 nsew
rlabel metal2 s 582166 -960 582278 480 4 la_oen[127]
port 432 nsew
rlabel metal2 s 171754 -960 171866 480 4 la_oen[12]
port 433 nsew
rlabel metal2 s 175342 -960 175454 480 4 la_oen[13]
port 434 nsew
rlabel metal2 s 178930 -960 179042 480 4 la_oen[14]
port 435 nsew
rlabel metal2 s 182518 -960 182630 480 4 la_oen[15]
port 436 nsew
rlabel metal2 s 186014 -960 186126 480 4 la_oen[16]
port 437 nsew
rlabel metal2 s 189602 -960 189714 480 4 la_oen[17]
port 438 nsew
rlabel metal2 s 193190 -960 193302 480 4 la_oen[18]
port 439 nsew
rlabel metal2 s 196778 -960 196890 480 4 la_oen[19]
port 440 nsew
rlabel metal2 s 132562 -960 132674 480 4 la_oen[1]
port 441 nsew
rlabel metal2 s 200366 -960 200478 480 4 la_oen[20]
port 442 nsew
rlabel metal2 s 203862 -960 203974 480 4 la_oen[21]
port 443 nsew
rlabel metal2 s 207450 -960 207562 480 4 la_oen[22]
port 444 nsew
rlabel metal2 s 211038 -960 211150 480 4 la_oen[23]
port 445 nsew
rlabel metal2 s 214626 -960 214738 480 4 la_oen[24]
port 446 nsew
rlabel metal2 s 218122 -960 218234 480 4 la_oen[25]
port 447 nsew
rlabel metal2 s 221710 -960 221822 480 4 la_oen[26]
port 448 nsew
rlabel metal2 s 225298 -960 225410 480 4 la_oen[27]
port 449 nsew
rlabel metal2 s 228886 -960 228998 480 4 la_oen[28]
port 450 nsew
rlabel metal2 s 232474 -960 232586 480 4 la_oen[29]
port 451 nsew
rlabel metal2 s 136058 -960 136170 480 4 la_oen[2]
port 452 nsew
rlabel metal2 s 235970 -960 236082 480 4 la_oen[30]
port 453 nsew
rlabel metal2 s 239558 -960 239670 480 4 la_oen[31]
port 454 nsew
rlabel metal2 s 243146 -960 243258 480 4 la_oen[32]
port 455 nsew
rlabel metal2 s 246734 -960 246846 480 4 la_oen[33]
port 456 nsew
rlabel metal2 s 250322 -960 250434 480 4 la_oen[34]
port 457 nsew
rlabel metal2 s 253818 -960 253930 480 4 la_oen[35]
port 458 nsew
rlabel metal2 s 257406 -960 257518 480 4 la_oen[36]
port 459 nsew
rlabel metal2 s 260994 -960 261106 480 4 la_oen[37]
port 460 nsew
rlabel metal2 s 264582 -960 264694 480 4 la_oen[38]
port 461 nsew
rlabel metal2 s 268078 -960 268190 480 4 la_oen[39]
port 462 nsew
rlabel metal2 s 139646 -960 139758 480 4 la_oen[3]
port 463 nsew
rlabel metal2 s 271666 -960 271778 480 4 la_oen[40]
port 464 nsew
rlabel metal2 s 275254 -960 275366 480 4 la_oen[41]
port 465 nsew
rlabel metal2 s 278842 -960 278954 480 4 la_oen[42]
port 466 nsew
rlabel metal2 s 282430 -960 282542 480 4 la_oen[43]
port 467 nsew
rlabel metal2 s 285926 -960 286038 480 4 la_oen[44]
port 468 nsew
rlabel metal2 s 289514 -960 289626 480 4 la_oen[45]
port 469 nsew
rlabel metal2 s 293102 -960 293214 480 4 la_oen[46]
port 470 nsew
rlabel metal2 s 296690 -960 296802 480 4 la_oen[47]
port 471 nsew
rlabel metal2 s 300278 -960 300390 480 4 la_oen[48]
port 472 nsew
rlabel metal2 s 303774 -960 303886 480 4 la_oen[49]
port 473 nsew
rlabel metal2 s 143234 -960 143346 480 4 la_oen[4]
port 474 nsew
rlabel metal2 s 307362 -960 307474 480 4 la_oen[50]
port 475 nsew
rlabel metal2 s 310950 -960 311062 480 4 la_oen[51]
port 476 nsew
rlabel metal2 s 314538 -960 314650 480 4 la_oen[52]
port 477 nsew
rlabel metal2 s 318034 -960 318146 480 4 la_oen[53]
port 478 nsew
rlabel metal2 s 321622 -960 321734 480 4 la_oen[54]
port 479 nsew
rlabel metal2 s 325210 -960 325322 480 4 la_oen[55]
port 480 nsew
rlabel metal2 s 328798 -960 328910 480 4 la_oen[56]
port 481 nsew
rlabel metal2 s 332386 -960 332498 480 4 la_oen[57]
port 482 nsew
rlabel metal2 s 335882 -960 335994 480 4 la_oen[58]
port 483 nsew
rlabel metal2 s 339470 -960 339582 480 4 la_oen[59]
port 484 nsew
rlabel metal2 s 146822 -960 146934 480 4 la_oen[5]
port 485 nsew
rlabel metal2 s 343058 -960 343170 480 4 la_oen[60]
port 486 nsew
rlabel metal2 s 346646 -960 346758 480 4 la_oen[61]
port 487 nsew
rlabel metal2 s 350234 -960 350346 480 4 la_oen[62]
port 488 nsew
rlabel metal2 s 353730 -960 353842 480 4 la_oen[63]
port 489 nsew
rlabel metal2 s 357318 -960 357430 480 4 la_oen[64]
port 490 nsew
rlabel metal2 s 360906 -960 361018 480 4 la_oen[65]
port 491 nsew
rlabel metal2 s 364494 -960 364606 480 4 la_oen[66]
port 492 nsew
rlabel metal2 s 367990 -960 368102 480 4 la_oen[67]
port 493 nsew
rlabel metal2 s 371578 -960 371690 480 4 la_oen[68]
port 494 nsew
rlabel metal2 s 375166 -960 375278 480 4 la_oen[69]
port 495 nsew
rlabel metal2 s 150410 -960 150522 480 4 la_oen[6]
port 496 nsew
rlabel metal2 s 378754 -960 378866 480 4 la_oen[70]
port 497 nsew
rlabel metal2 s 382342 -960 382454 480 4 la_oen[71]
port 498 nsew
rlabel metal2 s 385838 -960 385950 480 4 la_oen[72]
port 499 nsew
rlabel metal2 s 389426 -960 389538 480 4 la_oen[73]
port 500 nsew
rlabel metal2 s 393014 -960 393126 480 4 la_oen[74]
port 501 nsew
rlabel metal2 s 396602 -960 396714 480 4 la_oen[75]
port 502 nsew
rlabel metal2 s 400190 -960 400302 480 4 la_oen[76]
port 503 nsew
rlabel metal2 s 403686 -960 403798 480 4 la_oen[77]
port 504 nsew
rlabel metal2 s 407274 -960 407386 480 4 la_oen[78]
port 505 nsew
rlabel metal2 s 410862 -960 410974 480 4 la_oen[79]
port 506 nsew
rlabel metal2 s 153906 -960 154018 480 4 la_oen[7]
port 507 nsew
rlabel metal2 s 414450 -960 414562 480 4 la_oen[80]
port 508 nsew
rlabel metal2 s 417946 -960 418058 480 4 la_oen[81]
port 509 nsew
rlabel metal2 s 421534 -960 421646 480 4 la_oen[82]
port 510 nsew
rlabel metal2 s 425122 -960 425234 480 4 la_oen[83]
port 511 nsew
rlabel metal2 s 428710 -960 428822 480 4 la_oen[84]
port 512 nsew
rlabel metal2 s 432298 -960 432410 480 4 la_oen[85]
port 513 nsew
rlabel metal2 s 435794 -960 435906 480 4 la_oen[86]
port 514 nsew
rlabel metal2 s 439382 -960 439494 480 4 la_oen[87]
port 515 nsew
rlabel metal2 s 442970 -960 443082 480 4 la_oen[88]
port 516 nsew
rlabel metal2 s 446558 -960 446670 480 4 la_oen[89]
port 517 nsew
rlabel metal2 s 157494 -960 157606 480 4 la_oen[8]
port 518 nsew
rlabel metal2 s 450146 -960 450258 480 4 la_oen[90]
port 519 nsew
rlabel metal2 s 453642 -960 453754 480 4 la_oen[91]
port 520 nsew
rlabel metal2 s 457230 -960 457342 480 4 la_oen[92]
port 521 nsew
rlabel metal2 s 460818 -960 460930 480 4 la_oen[93]
port 522 nsew
rlabel metal2 s 464406 -960 464518 480 4 la_oen[94]
port 523 nsew
rlabel metal2 s 467902 -960 468014 480 4 la_oen[95]
port 524 nsew
rlabel metal2 s 471490 -960 471602 480 4 la_oen[96]
port 525 nsew
rlabel metal2 s 475078 -960 475190 480 4 la_oen[97]
port 526 nsew
rlabel metal2 s 478666 -960 478778 480 4 la_oen[98]
port 527 nsew
rlabel metal2 s 482254 -960 482366 480 4 la_oen[99]
port 528 nsew
rlabel metal2 s 161082 -960 161194 480 4 la_oen[9]
port 529 nsew
rlabel metal2 s 583362 -960 583474 480 4 user_clock2
port 530 nsew
rlabel metal2 s 542 -960 654 480 4 wb_clk_i
port 531 nsew
rlabel metal2 s 1646 -960 1758 480 4 wb_rst_i
port 532 nsew
rlabel metal2 s 2842 -960 2954 480 4 wbs_ack_o
port 533 nsew
rlabel metal2 s 7626 -960 7738 480 4 wbs_adr_i[0]
port 534 nsew
rlabel metal2 s 48106 -960 48218 480 4 wbs_adr_i[10]
port 535 nsew
rlabel metal2 s 51602 -960 51714 480 4 wbs_adr_i[11]
port 536 nsew
rlabel metal2 s 55190 -960 55302 480 4 wbs_adr_i[12]
port 537 nsew
rlabel metal2 s 58778 -960 58890 480 4 wbs_adr_i[13]
port 538 nsew
rlabel metal2 s 62366 -960 62478 480 4 wbs_adr_i[14]
port 539 nsew
rlabel metal2 s 65954 -960 66066 480 4 wbs_adr_i[15]
port 540 nsew
rlabel metal2 s 69450 -960 69562 480 4 wbs_adr_i[16]
port 541 nsew
rlabel metal2 s 73038 -960 73150 480 4 wbs_adr_i[17]
port 542 nsew
rlabel metal2 s 76626 -960 76738 480 4 wbs_adr_i[18]
port 543 nsew
rlabel metal2 s 80214 -960 80326 480 4 wbs_adr_i[19]
port 544 nsew
rlabel metal2 s 12410 -960 12522 480 4 wbs_adr_i[1]
port 545 nsew
rlabel metal2 s 83802 -960 83914 480 4 wbs_adr_i[20]
port 546 nsew
rlabel metal2 s 87298 -960 87410 480 4 wbs_adr_i[21]
port 547 nsew
rlabel metal2 s 90886 -960 90998 480 4 wbs_adr_i[22]
port 548 nsew
rlabel metal2 s 94474 -960 94586 480 4 wbs_adr_i[23]
port 549 nsew
rlabel metal2 s 98062 -960 98174 480 4 wbs_adr_i[24]
port 550 nsew
rlabel metal2 s 101558 -960 101670 480 4 wbs_adr_i[25]
port 551 nsew
rlabel metal2 s 105146 -960 105258 480 4 wbs_adr_i[26]
port 552 nsew
rlabel metal2 s 108734 -960 108846 480 4 wbs_adr_i[27]
port 553 nsew
rlabel metal2 s 112322 -960 112434 480 4 wbs_adr_i[28]
port 554 nsew
rlabel metal2 s 115910 -960 116022 480 4 wbs_adr_i[29]
port 555 nsew
rlabel metal2 s 17194 -960 17306 480 4 wbs_adr_i[2]
port 556 nsew
rlabel metal2 s 119406 -960 119518 480 4 wbs_adr_i[30]
port 557 nsew
rlabel metal2 s 122994 -960 123106 480 4 wbs_adr_i[31]
port 558 nsew
rlabel metal2 s 21886 -960 21998 480 4 wbs_adr_i[3]
port 559 nsew
rlabel metal2 s 26670 -960 26782 480 4 wbs_adr_i[4]
port 560 nsew
rlabel metal2 s 30258 -960 30370 480 4 wbs_adr_i[5]
port 561 nsew
rlabel metal2 s 33846 -960 33958 480 4 wbs_adr_i[6]
port 562 nsew
rlabel metal2 s 37342 -960 37454 480 4 wbs_adr_i[7]
port 563 nsew
rlabel metal2 s 40930 -960 41042 480 4 wbs_adr_i[8]
port 564 nsew
rlabel metal2 s 44518 -960 44630 480 4 wbs_adr_i[9]
port 565 nsew
rlabel metal2 s 4038 -960 4150 480 4 wbs_cyc_i
port 566 nsew
rlabel metal2 s 8822 -960 8934 480 4 wbs_dat_i[0]
port 567 nsew
rlabel metal2 s 49302 -960 49414 480 4 wbs_dat_i[10]
port 568 nsew
rlabel metal2 s 52798 -960 52910 480 4 wbs_dat_i[11]
port 569 nsew
rlabel metal2 s 56386 -960 56498 480 4 wbs_dat_i[12]
port 570 nsew
rlabel metal2 s 59974 -960 60086 480 4 wbs_dat_i[13]
port 571 nsew
rlabel metal2 s 63562 -960 63674 480 4 wbs_dat_i[14]
port 572 nsew
rlabel metal2 s 67150 -960 67262 480 4 wbs_dat_i[15]
port 573 nsew
rlabel metal2 s 70646 -960 70758 480 4 wbs_dat_i[16]
port 574 nsew
rlabel metal2 s 74234 -960 74346 480 4 wbs_dat_i[17]
port 575 nsew
rlabel metal2 s 77822 -960 77934 480 4 wbs_dat_i[18]
port 576 nsew
rlabel metal2 s 81410 -960 81522 480 4 wbs_dat_i[19]
port 577 nsew
rlabel metal2 s 13606 -960 13718 480 4 wbs_dat_i[1]
port 578 nsew
rlabel metal2 s 84906 -960 85018 480 4 wbs_dat_i[20]
port 579 nsew
rlabel metal2 s 88494 -960 88606 480 4 wbs_dat_i[21]
port 580 nsew
rlabel metal2 s 92082 -960 92194 480 4 wbs_dat_i[22]
port 581 nsew
rlabel metal2 s 95670 -960 95782 480 4 wbs_dat_i[23]
port 582 nsew
rlabel metal2 s 99258 -960 99370 480 4 wbs_dat_i[24]
port 583 nsew
rlabel metal2 s 102754 -960 102866 480 4 wbs_dat_i[25]
port 584 nsew
rlabel metal2 s 106342 -960 106454 480 4 wbs_dat_i[26]
port 585 nsew
rlabel metal2 s 109930 -960 110042 480 4 wbs_dat_i[27]
port 586 nsew
rlabel metal2 s 113518 -960 113630 480 4 wbs_dat_i[28]
port 587 nsew
rlabel metal2 s 117106 -960 117218 480 4 wbs_dat_i[29]
port 588 nsew
rlabel metal2 s 18298 -960 18410 480 4 wbs_dat_i[2]
port 589 nsew
rlabel metal2 s 120602 -960 120714 480 4 wbs_dat_i[30]
port 590 nsew
rlabel metal2 s 124190 -960 124302 480 4 wbs_dat_i[31]
port 591 nsew
rlabel metal2 s 23082 -960 23194 480 4 wbs_dat_i[3]
port 592 nsew
rlabel metal2 s 27866 -960 27978 480 4 wbs_dat_i[4]
port 593 nsew
rlabel metal2 s 31454 -960 31566 480 4 wbs_dat_i[5]
port 594 nsew
rlabel metal2 s 34950 -960 35062 480 4 wbs_dat_i[6]
port 595 nsew
rlabel metal2 s 38538 -960 38650 480 4 wbs_dat_i[7]
port 596 nsew
rlabel metal2 s 42126 -960 42238 480 4 wbs_dat_i[8]
port 597 nsew
rlabel metal2 s 45714 -960 45826 480 4 wbs_dat_i[9]
port 598 nsew
rlabel metal2 s 10018 -960 10130 480 4 wbs_dat_o[0]
port 599 nsew
rlabel metal2 s 50498 -960 50610 480 4 wbs_dat_o[10]
port 600 nsew
rlabel metal2 s 53994 -960 54106 480 4 wbs_dat_o[11]
port 601 nsew
rlabel metal2 s 57582 -960 57694 480 4 wbs_dat_o[12]
port 602 nsew
rlabel metal2 s 61170 -960 61282 480 4 wbs_dat_o[13]
port 603 nsew
rlabel metal2 s 64758 -960 64870 480 4 wbs_dat_o[14]
port 604 nsew
rlabel metal2 s 68254 -960 68366 480 4 wbs_dat_o[15]
port 605 nsew
rlabel metal2 s 71842 -960 71954 480 4 wbs_dat_o[16]
port 606 nsew
rlabel metal2 s 75430 -960 75542 480 4 wbs_dat_o[17]
port 607 nsew
rlabel metal2 s 79018 -960 79130 480 4 wbs_dat_o[18]
port 608 nsew
rlabel metal2 s 82606 -960 82718 480 4 wbs_dat_o[19]
port 609 nsew
rlabel metal2 s 14802 -960 14914 480 4 wbs_dat_o[1]
port 610 nsew
rlabel metal2 s 86102 -960 86214 480 4 wbs_dat_o[20]
port 611 nsew
rlabel metal2 s 89690 -960 89802 480 4 wbs_dat_o[21]
port 612 nsew
rlabel metal2 s 93278 -960 93390 480 4 wbs_dat_o[22]
port 613 nsew
rlabel metal2 s 96866 -960 96978 480 4 wbs_dat_o[23]
port 614 nsew
rlabel metal2 s 100454 -960 100566 480 4 wbs_dat_o[24]
port 615 nsew
rlabel metal2 s 103950 -960 104062 480 4 wbs_dat_o[25]
port 616 nsew
rlabel metal2 s 107538 -960 107650 480 4 wbs_dat_o[26]
port 617 nsew
rlabel metal2 s 111126 -960 111238 480 4 wbs_dat_o[27]
port 618 nsew
rlabel metal2 s 114714 -960 114826 480 4 wbs_dat_o[28]
port 619 nsew
rlabel metal2 s 118210 -960 118322 480 4 wbs_dat_o[29]
port 620 nsew
rlabel metal2 s 19494 -960 19606 480 4 wbs_dat_o[2]
port 621 nsew
rlabel metal2 s 121798 -960 121910 480 4 wbs_dat_o[30]
port 622 nsew
rlabel metal2 s 125386 -960 125498 480 4 wbs_dat_o[31]
port 623 nsew
rlabel metal2 s 24278 -960 24390 480 4 wbs_dat_o[3]
port 624 nsew
rlabel metal2 s 29062 -960 29174 480 4 wbs_dat_o[4]
port 625 nsew
rlabel metal2 s 32650 -960 32762 480 4 wbs_dat_o[5]
port 626 nsew
rlabel metal2 s 36146 -960 36258 480 4 wbs_dat_o[6]
port 627 nsew
rlabel metal2 s 39734 -960 39846 480 4 wbs_dat_o[7]
port 628 nsew
rlabel metal2 s 43322 -960 43434 480 4 wbs_dat_o[8]
port 629 nsew
rlabel metal2 s 46910 -960 47022 480 4 wbs_dat_o[9]
port 630 nsew
rlabel metal2 s 11214 -960 11326 480 4 wbs_sel_i[0]
port 631 nsew
rlabel metal2 s 15998 -960 16110 480 4 wbs_sel_i[1]
port 632 nsew
rlabel metal2 s 20690 -960 20802 480 4 wbs_sel_i[2]
port 633 nsew
rlabel metal2 s 25474 -960 25586 480 4 wbs_sel_i[3]
port 634 nsew
rlabel metal2 s 5234 -960 5346 480 4 wbs_stb_i
port 635 nsew
rlabel metal2 s 6430 -960 6542 480 4 wbs_we_i
port 636 nsew
rlabel metal5 s -1996 -924 585920 -324 4 vccd1
port 637 nsew
rlabel metal5 s -2916 -1844 586840 -1244 4 vssd1
port 638 nsew
rlabel metal5 s -3836 -2764 587760 -2164 4 vccd2
port 639 nsew
rlabel metal5 s -4756 -3684 588680 -3084 4 vssd2
port 640 nsew
rlabel metal5 s -5676 -4604 589600 -4004 4 vdda1
port 641 nsew
rlabel metal5 s -6596 -5524 590520 -4924 4 vssa1
port 642 nsew
rlabel metal5 s -7516 -6444 591440 -5844 4 vdda2
port 643 nsew
rlabel metal5 s -8436 -7364 592360 -6764 4 vssa2
port 644 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string GDS_FILE /project/openlane/user_project_wrapper/runs/user_project_wrapper/results/magic/user_project_wrapper.gds
string GDS_END 15349614
string GDS_START 12480028
<< end >>
