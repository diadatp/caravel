magic
tech sky130A
magscale 1 2
timestamp 1608124816
<< obsli1 >>
rect 998 2159 118758 117521
<< obsm1 >>
rect 0 892 119480 117552
<< metal2 >>
rect 372 119200 428 120000
rect 1384 119200 1440 120000
rect 2396 119200 2452 120000
rect 3500 119200 3556 120000
rect 4512 119200 4568 120000
rect 5616 119200 5672 120000
rect 6628 119200 6684 120000
rect 7732 119200 7788 120000
rect 8744 119200 8800 120000
rect 9756 119200 9812 120000
rect 10860 119200 10916 120000
rect 11872 119200 11928 120000
rect 12976 119200 13032 120000
rect 13988 119200 14044 120000
rect 15092 119200 15148 120000
rect 16104 119200 16160 120000
rect 17208 119200 17264 120000
rect 18220 119200 18276 120000
rect 19232 119200 19288 120000
rect 20336 119200 20392 120000
rect 21348 119200 21404 120000
rect 22452 119200 22508 120000
rect 23464 119200 23520 120000
rect 24568 119200 24624 120000
rect 25580 119200 25636 120000
rect 26592 119200 26648 120000
rect 27696 119200 27752 120000
rect 28708 119200 28764 120000
rect 29812 119200 29868 120000
rect 30824 119200 30880 120000
rect 31928 119200 31984 120000
rect 32940 119200 32996 120000
rect 34044 119200 34100 120000
rect 35056 119200 35112 120000
rect 36068 119200 36124 120000
rect 37172 119200 37228 120000
rect 38184 119200 38240 120000
rect 39288 119200 39344 120000
rect 40300 119200 40356 120000
rect 41404 119200 41460 120000
rect 42416 119200 42472 120000
rect 43428 119200 43484 120000
rect 44532 119200 44588 120000
rect 45544 119200 45600 120000
rect 46648 119200 46704 120000
rect 47660 119200 47716 120000
rect 48764 119200 48820 120000
rect 49776 119200 49832 120000
rect 50880 119200 50936 120000
rect 51892 119200 51948 120000
rect 52904 119200 52960 120000
rect 54008 119200 54064 120000
rect 55020 119200 55076 120000
rect 56124 119200 56180 120000
rect 57136 119200 57192 120000
rect 58240 119200 58296 120000
rect 59252 119200 59308 120000
rect 60356 119200 60412 120000
rect 61368 119200 61424 120000
rect 62380 119200 62436 120000
rect 63484 119200 63540 120000
rect 64496 119200 64552 120000
rect 65600 119200 65656 120000
rect 66612 119200 66668 120000
rect 67716 119200 67772 120000
rect 68728 119200 68784 120000
rect 69740 119200 69796 120000
rect 70844 119200 70900 120000
rect 71856 119200 71912 120000
rect 72960 119200 73016 120000
rect 73972 119200 74028 120000
rect 75076 119200 75132 120000
rect 76088 119200 76144 120000
rect 77192 119200 77248 120000
rect 78204 119200 78260 120000
rect 79216 119200 79272 120000
rect 80320 119200 80376 120000
rect 81332 119200 81388 120000
rect 82436 119200 82492 120000
rect 83448 119200 83504 120000
rect 84552 119200 84608 120000
rect 85564 119200 85620 120000
rect 86576 119200 86632 120000
rect 87680 119200 87736 120000
rect 88692 119200 88748 120000
rect 89796 119200 89852 120000
rect 90808 119200 90864 120000
rect 91912 119200 91968 120000
rect 92924 119200 92980 120000
rect 94028 119200 94084 120000
rect 95040 119200 95096 120000
rect 96052 119200 96108 120000
rect 97156 119200 97212 120000
rect 98168 119200 98224 120000
rect 99272 119200 99328 120000
rect 100284 119200 100340 120000
rect 101388 119200 101444 120000
rect 102400 119200 102456 120000
rect 103412 119200 103468 120000
rect 104516 119200 104572 120000
rect 105528 119200 105584 120000
rect 106632 119200 106688 120000
rect 107644 119200 107700 120000
rect 108748 119200 108804 120000
rect 109760 119200 109816 120000
rect 110864 119200 110920 120000
rect 111876 119200 111932 120000
rect 112888 119200 112944 120000
rect 113992 119200 114048 120000
rect 115004 119200 115060 120000
rect 116108 119200 116164 120000
rect 117120 119200 117176 120000
rect 118224 119200 118280 120000
rect 119236 119200 119292 120000
rect 4 0 60 800
rect 188 0 244 800
rect 464 0 520 800
rect 648 0 704 800
rect 924 0 980 800
rect 1200 0 1256 800
rect 1384 0 1440 800
rect 1660 0 1716 800
rect 1936 0 1992 800
rect 2120 0 2176 800
rect 2396 0 2452 800
rect 2672 0 2728 800
rect 2856 0 2912 800
rect 3132 0 3188 800
rect 3408 0 3464 800
rect 3592 0 3648 800
rect 3868 0 3924 800
rect 4144 0 4200 800
rect 4328 0 4384 800
rect 4604 0 4660 800
rect 4880 0 4936 800
rect 5064 0 5120 800
rect 5340 0 5396 800
rect 5616 0 5672 800
rect 5800 0 5856 800
rect 6076 0 6132 800
rect 6352 0 6408 800
rect 6536 0 6592 800
rect 6812 0 6868 800
rect 7088 0 7144 800
rect 7272 0 7328 800
rect 7548 0 7604 800
rect 7824 0 7880 800
rect 8008 0 8064 800
rect 8284 0 8340 800
rect 8560 0 8616 800
rect 8744 0 8800 800
rect 9020 0 9076 800
rect 9296 0 9352 800
rect 9480 0 9536 800
rect 9756 0 9812 800
rect 10032 0 10088 800
rect 10216 0 10272 800
rect 10492 0 10548 800
rect 10768 0 10824 800
rect 10952 0 11008 800
rect 11228 0 11284 800
rect 11504 0 11560 800
rect 11688 0 11744 800
rect 11964 0 12020 800
rect 12240 0 12296 800
rect 12424 0 12480 800
rect 12700 0 12756 800
rect 12976 0 13032 800
rect 13160 0 13216 800
rect 13436 0 13492 800
rect 13712 0 13768 800
rect 13896 0 13952 800
rect 14172 0 14228 800
rect 14448 0 14504 800
rect 14632 0 14688 800
rect 14908 0 14964 800
rect 15092 0 15148 800
rect 15368 0 15424 800
rect 15644 0 15700 800
rect 15828 0 15884 800
rect 16104 0 16160 800
rect 16380 0 16436 800
rect 16564 0 16620 800
rect 16840 0 16896 800
rect 17116 0 17172 800
rect 17300 0 17356 800
rect 17576 0 17632 800
rect 17852 0 17908 800
rect 18036 0 18092 800
rect 18312 0 18368 800
rect 18588 0 18644 800
rect 18772 0 18828 800
rect 19048 0 19104 800
rect 19324 0 19380 800
rect 19508 0 19564 800
rect 19784 0 19840 800
rect 20060 0 20116 800
rect 20244 0 20300 800
rect 20520 0 20576 800
rect 20796 0 20852 800
rect 20980 0 21036 800
rect 21256 0 21312 800
rect 21532 0 21588 800
rect 21716 0 21772 800
rect 21992 0 22048 800
rect 22268 0 22324 800
rect 22452 0 22508 800
rect 22728 0 22784 800
rect 23004 0 23060 800
rect 23188 0 23244 800
rect 23464 0 23520 800
rect 23740 0 23796 800
rect 23924 0 23980 800
rect 24200 0 24256 800
rect 24476 0 24532 800
rect 24660 0 24716 800
rect 24936 0 24992 800
rect 25212 0 25268 800
rect 25396 0 25452 800
rect 25672 0 25728 800
rect 25948 0 26004 800
rect 26132 0 26188 800
rect 26408 0 26464 800
rect 26684 0 26740 800
rect 26868 0 26924 800
rect 27144 0 27200 800
rect 27420 0 27476 800
rect 27604 0 27660 800
rect 27880 0 27936 800
rect 28156 0 28212 800
rect 28340 0 28396 800
rect 28616 0 28672 800
rect 28892 0 28948 800
rect 29076 0 29132 800
rect 29352 0 29408 800
rect 29628 0 29684 800
rect 29812 0 29868 800
rect 30088 0 30144 800
rect 30272 0 30328 800
rect 30548 0 30604 800
rect 30824 0 30880 800
rect 31008 0 31064 800
rect 31284 0 31340 800
rect 31560 0 31616 800
rect 31744 0 31800 800
rect 32020 0 32076 800
rect 32296 0 32352 800
rect 32480 0 32536 800
rect 32756 0 32812 800
rect 33032 0 33088 800
rect 33216 0 33272 800
rect 33492 0 33548 800
rect 33768 0 33824 800
rect 33952 0 34008 800
rect 34228 0 34284 800
rect 34504 0 34560 800
rect 34688 0 34744 800
rect 34964 0 35020 800
rect 35240 0 35296 800
rect 35424 0 35480 800
rect 35700 0 35756 800
rect 35976 0 36032 800
rect 36160 0 36216 800
rect 36436 0 36492 800
rect 36712 0 36768 800
rect 36896 0 36952 800
rect 37172 0 37228 800
rect 37448 0 37504 800
rect 37632 0 37688 800
rect 37908 0 37964 800
rect 38184 0 38240 800
rect 38368 0 38424 800
rect 38644 0 38700 800
rect 38920 0 38976 800
rect 39104 0 39160 800
rect 39380 0 39436 800
rect 39656 0 39712 800
rect 39840 0 39896 800
rect 40116 0 40172 800
rect 40392 0 40448 800
rect 40576 0 40632 800
rect 40852 0 40908 800
rect 41128 0 41184 800
rect 41312 0 41368 800
rect 41588 0 41644 800
rect 41864 0 41920 800
rect 42048 0 42104 800
rect 42324 0 42380 800
rect 42600 0 42656 800
rect 42784 0 42840 800
rect 43060 0 43116 800
rect 43336 0 43392 800
rect 43520 0 43576 800
rect 43796 0 43852 800
rect 44072 0 44128 800
rect 44256 0 44312 800
rect 44532 0 44588 800
rect 44808 0 44864 800
rect 44992 0 45048 800
rect 45268 0 45324 800
rect 45452 0 45508 800
rect 45728 0 45784 800
rect 46004 0 46060 800
rect 46188 0 46244 800
rect 46464 0 46520 800
rect 46740 0 46796 800
rect 46924 0 46980 800
rect 47200 0 47256 800
rect 47476 0 47532 800
rect 47660 0 47716 800
rect 47936 0 47992 800
rect 48212 0 48268 800
rect 48396 0 48452 800
rect 48672 0 48728 800
rect 48948 0 49004 800
rect 49132 0 49188 800
rect 49408 0 49464 800
rect 49684 0 49740 800
rect 49868 0 49924 800
rect 50144 0 50200 800
rect 50420 0 50476 800
rect 50604 0 50660 800
rect 50880 0 50936 800
rect 51156 0 51212 800
rect 51340 0 51396 800
rect 51616 0 51672 800
rect 51892 0 51948 800
rect 52076 0 52132 800
rect 52352 0 52408 800
rect 52628 0 52684 800
rect 52812 0 52868 800
rect 53088 0 53144 800
rect 53364 0 53420 800
rect 53548 0 53604 800
rect 53824 0 53880 800
rect 54100 0 54156 800
rect 54284 0 54340 800
rect 54560 0 54616 800
rect 54836 0 54892 800
rect 55020 0 55076 800
rect 55296 0 55352 800
rect 55572 0 55628 800
rect 55756 0 55812 800
rect 56032 0 56088 800
rect 56308 0 56364 800
rect 56492 0 56548 800
rect 56768 0 56824 800
rect 57044 0 57100 800
rect 57228 0 57284 800
rect 57504 0 57560 800
rect 57780 0 57836 800
rect 57964 0 58020 800
rect 58240 0 58296 800
rect 58516 0 58572 800
rect 58700 0 58756 800
rect 58976 0 59032 800
rect 59252 0 59308 800
rect 59436 0 59492 800
rect 59712 0 59768 800
rect 59988 0 60044 800
rect 60172 0 60228 800
rect 60448 0 60504 800
rect 60632 0 60688 800
rect 60908 0 60964 800
rect 61184 0 61240 800
rect 61368 0 61424 800
rect 61644 0 61700 800
rect 61920 0 61976 800
rect 62104 0 62160 800
rect 62380 0 62436 800
rect 62656 0 62712 800
rect 62840 0 62896 800
rect 63116 0 63172 800
rect 63392 0 63448 800
rect 63576 0 63632 800
rect 63852 0 63908 800
rect 64128 0 64184 800
rect 64312 0 64368 800
rect 64588 0 64644 800
rect 64864 0 64920 800
rect 65048 0 65104 800
rect 65324 0 65380 800
rect 65600 0 65656 800
rect 65784 0 65840 800
rect 66060 0 66116 800
rect 66336 0 66392 800
rect 66520 0 66576 800
rect 66796 0 66852 800
rect 67072 0 67128 800
rect 67256 0 67312 800
rect 67532 0 67588 800
rect 67808 0 67864 800
rect 67992 0 68048 800
rect 68268 0 68324 800
rect 68544 0 68600 800
rect 68728 0 68784 800
rect 69004 0 69060 800
rect 69280 0 69336 800
rect 69464 0 69520 800
rect 69740 0 69796 800
rect 70016 0 70072 800
rect 70200 0 70256 800
rect 70476 0 70532 800
rect 70752 0 70808 800
rect 70936 0 70992 800
rect 71212 0 71268 800
rect 71488 0 71544 800
rect 71672 0 71728 800
rect 71948 0 72004 800
rect 72224 0 72280 800
rect 72408 0 72464 800
rect 72684 0 72740 800
rect 72960 0 73016 800
rect 73144 0 73200 800
rect 73420 0 73476 800
rect 73696 0 73752 800
rect 73880 0 73936 800
rect 74156 0 74212 800
rect 74432 0 74488 800
rect 74616 0 74672 800
rect 74892 0 74948 800
rect 75076 0 75132 800
rect 75352 0 75408 800
rect 75628 0 75684 800
rect 75812 0 75868 800
rect 76088 0 76144 800
rect 76364 0 76420 800
rect 76548 0 76604 800
rect 76824 0 76880 800
rect 77100 0 77156 800
rect 77284 0 77340 800
rect 77560 0 77616 800
rect 77836 0 77892 800
rect 78020 0 78076 800
rect 78296 0 78352 800
rect 78572 0 78628 800
rect 78756 0 78812 800
rect 79032 0 79088 800
rect 79308 0 79364 800
rect 79492 0 79548 800
rect 79768 0 79824 800
rect 80044 0 80100 800
rect 80228 0 80284 800
rect 80504 0 80560 800
rect 80780 0 80836 800
rect 80964 0 81020 800
rect 81240 0 81296 800
rect 81516 0 81572 800
rect 81700 0 81756 800
rect 81976 0 82032 800
rect 82252 0 82308 800
rect 82436 0 82492 800
rect 82712 0 82768 800
rect 82988 0 83044 800
rect 83172 0 83228 800
rect 83448 0 83504 800
rect 83724 0 83780 800
rect 83908 0 83964 800
rect 84184 0 84240 800
rect 84460 0 84516 800
rect 84644 0 84700 800
rect 84920 0 84976 800
rect 85196 0 85252 800
rect 85380 0 85436 800
rect 85656 0 85712 800
rect 85932 0 85988 800
rect 86116 0 86172 800
rect 86392 0 86448 800
rect 86668 0 86724 800
rect 86852 0 86908 800
rect 87128 0 87184 800
rect 87404 0 87460 800
rect 87588 0 87644 800
rect 87864 0 87920 800
rect 88140 0 88196 800
rect 88324 0 88380 800
rect 88600 0 88656 800
rect 88876 0 88932 800
rect 89060 0 89116 800
rect 89336 0 89392 800
rect 89612 0 89668 800
rect 89796 0 89852 800
rect 90072 0 90128 800
rect 90256 0 90312 800
rect 90532 0 90588 800
rect 90808 0 90864 800
rect 90992 0 91048 800
rect 91268 0 91324 800
rect 91544 0 91600 800
rect 91728 0 91784 800
rect 92004 0 92060 800
rect 92280 0 92336 800
rect 92464 0 92520 800
rect 92740 0 92796 800
rect 93016 0 93072 800
rect 93200 0 93256 800
rect 93476 0 93532 800
rect 93752 0 93808 800
rect 93936 0 93992 800
rect 94212 0 94268 800
rect 94488 0 94544 800
rect 94672 0 94728 800
rect 94948 0 95004 800
rect 95224 0 95280 800
rect 95408 0 95464 800
rect 95684 0 95740 800
rect 95960 0 96016 800
rect 96144 0 96200 800
rect 96420 0 96476 800
rect 96696 0 96752 800
rect 96880 0 96936 800
rect 97156 0 97212 800
rect 97432 0 97488 800
rect 97616 0 97672 800
rect 97892 0 97948 800
rect 98168 0 98224 800
rect 98352 0 98408 800
rect 98628 0 98684 800
rect 98904 0 98960 800
rect 99088 0 99144 800
rect 99364 0 99420 800
rect 99640 0 99696 800
rect 99824 0 99880 800
rect 100100 0 100156 800
rect 100376 0 100432 800
rect 100560 0 100616 800
rect 100836 0 100892 800
rect 101112 0 101168 800
rect 101296 0 101352 800
rect 101572 0 101628 800
rect 101848 0 101904 800
rect 102032 0 102088 800
rect 102308 0 102364 800
rect 102584 0 102640 800
rect 102768 0 102824 800
rect 103044 0 103100 800
rect 103320 0 103376 800
rect 103504 0 103560 800
rect 103780 0 103836 800
rect 104056 0 104112 800
rect 104240 0 104296 800
rect 104516 0 104572 800
rect 104792 0 104848 800
rect 104976 0 105032 800
rect 105252 0 105308 800
rect 105436 0 105492 800
rect 105712 0 105768 800
rect 105988 0 106044 800
rect 106172 0 106228 800
rect 106448 0 106504 800
rect 106724 0 106780 800
rect 106908 0 106964 800
rect 107184 0 107240 800
rect 107460 0 107516 800
rect 107644 0 107700 800
rect 107920 0 107976 800
rect 108196 0 108252 800
rect 108380 0 108436 800
rect 108656 0 108712 800
rect 108932 0 108988 800
rect 109116 0 109172 800
rect 109392 0 109448 800
rect 109668 0 109724 800
rect 109852 0 109908 800
rect 110128 0 110184 800
rect 110404 0 110460 800
rect 110588 0 110644 800
rect 110864 0 110920 800
rect 111140 0 111196 800
rect 111324 0 111380 800
rect 111600 0 111656 800
rect 111876 0 111932 800
rect 112060 0 112116 800
rect 112336 0 112392 800
rect 112612 0 112668 800
rect 112796 0 112852 800
rect 113072 0 113128 800
rect 113348 0 113404 800
rect 113532 0 113588 800
rect 113808 0 113864 800
rect 114084 0 114140 800
rect 114268 0 114324 800
rect 114544 0 114600 800
rect 114820 0 114876 800
rect 115004 0 115060 800
rect 115280 0 115336 800
rect 115556 0 115612 800
rect 115740 0 115796 800
rect 116016 0 116072 800
rect 116292 0 116348 800
rect 116476 0 116532 800
rect 116752 0 116808 800
rect 117028 0 117084 800
rect 117212 0 117268 800
rect 117488 0 117544 800
rect 117764 0 117820 800
rect 117948 0 118004 800
rect 118224 0 118280 800
rect 118500 0 118556 800
rect 118684 0 118740 800
rect 118960 0 119016 800
rect 119236 0 119292 800
rect 119420 0 119476 800
rect 119696 0 119752 800
<< obsm2 >>
rect 6 119144 316 119200
rect 484 119144 1328 119200
rect 1496 119144 2340 119200
rect 2508 119144 3444 119200
rect 3612 119144 4456 119200
rect 4624 119144 5560 119200
rect 5728 119144 6572 119200
rect 6740 119144 7676 119200
rect 7844 119144 8688 119200
rect 8856 119144 9700 119200
rect 9868 119144 10804 119200
rect 10972 119144 11816 119200
rect 11984 119144 12920 119200
rect 13088 119144 13932 119200
rect 14100 119144 15036 119200
rect 15204 119144 16048 119200
rect 16216 119144 17152 119200
rect 17320 119144 18164 119200
rect 18332 119144 19176 119200
rect 19344 119144 20280 119200
rect 20448 119144 21292 119200
rect 21460 119144 22396 119200
rect 22564 119144 23408 119200
rect 23576 119144 24512 119200
rect 24680 119144 25524 119200
rect 25692 119144 26536 119200
rect 26704 119144 27640 119200
rect 27808 119144 28652 119200
rect 28820 119144 29756 119200
rect 29924 119144 30768 119200
rect 30936 119144 31872 119200
rect 32040 119144 32884 119200
rect 33052 119144 33988 119200
rect 34156 119144 35000 119200
rect 35168 119144 36012 119200
rect 36180 119144 37116 119200
rect 37284 119144 38128 119200
rect 38296 119144 39232 119200
rect 39400 119144 40244 119200
rect 40412 119144 41348 119200
rect 41516 119144 42360 119200
rect 42528 119144 43372 119200
rect 43540 119144 44476 119200
rect 44644 119144 45488 119200
rect 45656 119144 46592 119200
rect 46760 119144 47604 119200
rect 47772 119144 48708 119200
rect 48876 119144 49720 119200
rect 49888 119144 50824 119200
rect 50992 119144 51836 119200
rect 52004 119144 52848 119200
rect 53016 119144 53952 119200
rect 54120 119144 54964 119200
rect 55132 119144 56068 119200
rect 56236 119144 57080 119200
rect 57248 119144 58184 119200
rect 58352 119144 59196 119200
rect 59364 119144 60300 119200
rect 60468 119144 61312 119200
rect 61480 119144 62324 119200
rect 62492 119144 63428 119200
rect 63596 119144 64440 119200
rect 64608 119144 65544 119200
rect 65712 119144 66556 119200
rect 66724 119144 67660 119200
rect 67828 119144 68672 119200
rect 68840 119144 69684 119200
rect 69852 119144 70788 119200
rect 70956 119144 71800 119200
rect 71968 119144 72904 119200
rect 73072 119144 73916 119200
rect 74084 119144 75020 119200
rect 75188 119144 76032 119200
rect 76200 119144 77136 119200
rect 77304 119144 78148 119200
rect 78316 119144 79160 119200
rect 79328 119144 80264 119200
rect 80432 119144 81276 119200
rect 81444 119144 82380 119200
rect 82548 119144 83392 119200
rect 83560 119144 84496 119200
rect 84664 119144 85508 119200
rect 85676 119144 86520 119200
rect 86688 119144 87624 119200
rect 87792 119144 88636 119200
rect 88804 119144 89740 119200
rect 89908 119144 90752 119200
rect 90920 119144 91856 119200
rect 92024 119144 92868 119200
rect 93036 119144 93972 119200
rect 94140 119144 94984 119200
rect 95152 119144 95996 119200
rect 96164 119144 97100 119200
rect 97268 119144 98112 119200
rect 98280 119144 99216 119200
rect 99384 119144 100228 119200
rect 100396 119144 101332 119200
rect 101500 119144 102344 119200
rect 102512 119144 103356 119200
rect 103524 119144 104460 119200
rect 104628 119144 105472 119200
rect 105640 119144 106576 119200
rect 106744 119144 107588 119200
rect 107756 119144 108692 119200
rect 108860 119144 109704 119200
rect 109872 119144 110808 119200
rect 110976 119144 111820 119200
rect 111988 119144 112832 119200
rect 113000 119144 113936 119200
rect 114104 119144 114948 119200
rect 115116 119144 116052 119200
rect 116220 119144 117064 119200
rect 117232 119144 118168 119200
rect 118336 119144 119180 119200
rect 119348 119144 119474 119200
rect 6 856 119474 119144
rect 116 800 132 856
rect 300 800 408 856
rect 576 800 592 856
rect 760 800 868 856
rect 1036 800 1144 856
rect 1312 800 1328 856
rect 1496 800 1604 856
rect 1772 800 1880 856
rect 2048 800 2064 856
rect 2232 800 2340 856
rect 2508 800 2616 856
rect 2784 800 2800 856
rect 2968 800 3076 856
rect 3244 800 3352 856
rect 3520 800 3536 856
rect 3704 800 3812 856
rect 3980 800 4088 856
rect 4256 800 4272 856
rect 4440 800 4548 856
rect 4716 800 4824 856
rect 4992 800 5008 856
rect 5176 800 5284 856
rect 5452 800 5560 856
rect 5728 800 5744 856
rect 5912 800 6020 856
rect 6188 800 6296 856
rect 6464 800 6480 856
rect 6648 800 6756 856
rect 6924 800 7032 856
rect 7200 800 7216 856
rect 7384 800 7492 856
rect 7660 800 7768 856
rect 7936 800 7952 856
rect 8120 800 8228 856
rect 8396 800 8504 856
rect 8672 800 8688 856
rect 8856 800 8964 856
rect 9132 800 9240 856
rect 9408 800 9424 856
rect 9592 800 9700 856
rect 9868 800 9976 856
rect 10144 800 10160 856
rect 10328 800 10436 856
rect 10604 800 10712 856
rect 10880 800 10896 856
rect 11064 800 11172 856
rect 11340 800 11448 856
rect 11616 800 11632 856
rect 11800 800 11908 856
rect 12076 800 12184 856
rect 12352 800 12368 856
rect 12536 800 12644 856
rect 12812 800 12920 856
rect 13088 800 13104 856
rect 13272 800 13380 856
rect 13548 800 13656 856
rect 13824 800 13840 856
rect 14008 800 14116 856
rect 14284 800 14392 856
rect 14560 800 14576 856
rect 14744 800 14852 856
rect 15020 800 15036 856
rect 15204 800 15312 856
rect 15480 800 15588 856
rect 15756 800 15772 856
rect 15940 800 16048 856
rect 16216 800 16324 856
rect 16492 800 16508 856
rect 16676 800 16784 856
rect 16952 800 17060 856
rect 17228 800 17244 856
rect 17412 800 17520 856
rect 17688 800 17796 856
rect 17964 800 17980 856
rect 18148 800 18256 856
rect 18424 800 18532 856
rect 18700 800 18716 856
rect 18884 800 18992 856
rect 19160 800 19268 856
rect 19436 800 19452 856
rect 19620 800 19728 856
rect 19896 800 20004 856
rect 20172 800 20188 856
rect 20356 800 20464 856
rect 20632 800 20740 856
rect 20908 800 20924 856
rect 21092 800 21200 856
rect 21368 800 21476 856
rect 21644 800 21660 856
rect 21828 800 21936 856
rect 22104 800 22212 856
rect 22380 800 22396 856
rect 22564 800 22672 856
rect 22840 800 22948 856
rect 23116 800 23132 856
rect 23300 800 23408 856
rect 23576 800 23684 856
rect 23852 800 23868 856
rect 24036 800 24144 856
rect 24312 800 24420 856
rect 24588 800 24604 856
rect 24772 800 24880 856
rect 25048 800 25156 856
rect 25324 800 25340 856
rect 25508 800 25616 856
rect 25784 800 25892 856
rect 26060 800 26076 856
rect 26244 800 26352 856
rect 26520 800 26628 856
rect 26796 800 26812 856
rect 26980 800 27088 856
rect 27256 800 27364 856
rect 27532 800 27548 856
rect 27716 800 27824 856
rect 27992 800 28100 856
rect 28268 800 28284 856
rect 28452 800 28560 856
rect 28728 800 28836 856
rect 29004 800 29020 856
rect 29188 800 29296 856
rect 29464 800 29572 856
rect 29740 800 29756 856
rect 29924 800 30032 856
rect 30200 800 30216 856
rect 30384 800 30492 856
rect 30660 800 30768 856
rect 30936 800 30952 856
rect 31120 800 31228 856
rect 31396 800 31504 856
rect 31672 800 31688 856
rect 31856 800 31964 856
rect 32132 800 32240 856
rect 32408 800 32424 856
rect 32592 800 32700 856
rect 32868 800 32976 856
rect 33144 800 33160 856
rect 33328 800 33436 856
rect 33604 800 33712 856
rect 33880 800 33896 856
rect 34064 800 34172 856
rect 34340 800 34448 856
rect 34616 800 34632 856
rect 34800 800 34908 856
rect 35076 800 35184 856
rect 35352 800 35368 856
rect 35536 800 35644 856
rect 35812 800 35920 856
rect 36088 800 36104 856
rect 36272 800 36380 856
rect 36548 800 36656 856
rect 36824 800 36840 856
rect 37008 800 37116 856
rect 37284 800 37392 856
rect 37560 800 37576 856
rect 37744 800 37852 856
rect 38020 800 38128 856
rect 38296 800 38312 856
rect 38480 800 38588 856
rect 38756 800 38864 856
rect 39032 800 39048 856
rect 39216 800 39324 856
rect 39492 800 39600 856
rect 39768 800 39784 856
rect 39952 800 40060 856
rect 40228 800 40336 856
rect 40504 800 40520 856
rect 40688 800 40796 856
rect 40964 800 41072 856
rect 41240 800 41256 856
rect 41424 800 41532 856
rect 41700 800 41808 856
rect 41976 800 41992 856
rect 42160 800 42268 856
rect 42436 800 42544 856
rect 42712 800 42728 856
rect 42896 800 43004 856
rect 43172 800 43280 856
rect 43448 800 43464 856
rect 43632 800 43740 856
rect 43908 800 44016 856
rect 44184 800 44200 856
rect 44368 800 44476 856
rect 44644 800 44752 856
rect 44920 800 44936 856
rect 45104 800 45212 856
rect 45380 800 45396 856
rect 45564 800 45672 856
rect 45840 800 45948 856
rect 46116 800 46132 856
rect 46300 800 46408 856
rect 46576 800 46684 856
rect 46852 800 46868 856
rect 47036 800 47144 856
rect 47312 800 47420 856
rect 47588 800 47604 856
rect 47772 800 47880 856
rect 48048 800 48156 856
rect 48324 800 48340 856
rect 48508 800 48616 856
rect 48784 800 48892 856
rect 49060 800 49076 856
rect 49244 800 49352 856
rect 49520 800 49628 856
rect 49796 800 49812 856
rect 49980 800 50088 856
rect 50256 800 50364 856
rect 50532 800 50548 856
rect 50716 800 50824 856
rect 50992 800 51100 856
rect 51268 800 51284 856
rect 51452 800 51560 856
rect 51728 800 51836 856
rect 52004 800 52020 856
rect 52188 800 52296 856
rect 52464 800 52572 856
rect 52740 800 52756 856
rect 52924 800 53032 856
rect 53200 800 53308 856
rect 53476 800 53492 856
rect 53660 800 53768 856
rect 53936 800 54044 856
rect 54212 800 54228 856
rect 54396 800 54504 856
rect 54672 800 54780 856
rect 54948 800 54964 856
rect 55132 800 55240 856
rect 55408 800 55516 856
rect 55684 800 55700 856
rect 55868 800 55976 856
rect 56144 800 56252 856
rect 56420 800 56436 856
rect 56604 800 56712 856
rect 56880 800 56988 856
rect 57156 800 57172 856
rect 57340 800 57448 856
rect 57616 800 57724 856
rect 57892 800 57908 856
rect 58076 800 58184 856
rect 58352 800 58460 856
rect 58628 800 58644 856
rect 58812 800 58920 856
rect 59088 800 59196 856
rect 59364 800 59380 856
rect 59548 800 59656 856
rect 59824 800 59932 856
rect 60100 800 60116 856
rect 60284 800 60392 856
rect 60560 800 60576 856
rect 60744 800 60852 856
rect 61020 800 61128 856
rect 61296 800 61312 856
rect 61480 800 61588 856
rect 61756 800 61864 856
rect 62032 800 62048 856
rect 62216 800 62324 856
rect 62492 800 62600 856
rect 62768 800 62784 856
rect 62952 800 63060 856
rect 63228 800 63336 856
rect 63504 800 63520 856
rect 63688 800 63796 856
rect 63964 800 64072 856
rect 64240 800 64256 856
rect 64424 800 64532 856
rect 64700 800 64808 856
rect 64976 800 64992 856
rect 65160 800 65268 856
rect 65436 800 65544 856
rect 65712 800 65728 856
rect 65896 800 66004 856
rect 66172 800 66280 856
rect 66448 800 66464 856
rect 66632 800 66740 856
rect 66908 800 67016 856
rect 67184 800 67200 856
rect 67368 800 67476 856
rect 67644 800 67752 856
rect 67920 800 67936 856
rect 68104 800 68212 856
rect 68380 800 68488 856
rect 68656 800 68672 856
rect 68840 800 68948 856
rect 69116 800 69224 856
rect 69392 800 69408 856
rect 69576 800 69684 856
rect 69852 800 69960 856
rect 70128 800 70144 856
rect 70312 800 70420 856
rect 70588 800 70696 856
rect 70864 800 70880 856
rect 71048 800 71156 856
rect 71324 800 71432 856
rect 71600 800 71616 856
rect 71784 800 71892 856
rect 72060 800 72168 856
rect 72336 800 72352 856
rect 72520 800 72628 856
rect 72796 800 72904 856
rect 73072 800 73088 856
rect 73256 800 73364 856
rect 73532 800 73640 856
rect 73808 800 73824 856
rect 73992 800 74100 856
rect 74268 800 74376 856
rect 74544 800 74560 856
rect 74728 800 74836 856
rect 75004 800 75020 856
rect 75188 800 75296 856
rect 75464 800 75572 856
rect 75740 800 75756 856
rect 75924 800 76032 856
rect 76200 800 76308 856
rect 76476 800 76492 856
rect 76660 800 76768 856
rect 76936 800 77044 856
rect 77212 800 77228 856
rect 77396 800 77504 856
rect 77672 800 77780 856
rect 77948 800 77964 856
rect 78132 800 78240 856
rect 78408 800 78516 856
rect 78684 800 78700 856
rect 78868 800 78976 856
rect 79144 800 79252 856
rect 79420 800 79436 856
rect 79604 800 79712 856
rect 79880 800 79988 856
rect 80156 800 80172 856
rect 80340 800 80448 856
rect 80616 800 80724 856
rect 80892 800 80908 856
rect 81076 800 81184 856
rect 81352 800 81460 856
rect 81628 800 81644 856
rect 81812 800 81920 856
rect 82088 800 82196 856
rect 82364 800 82380 856
rect 82548 800 82656 856
rect 82824 800 82932 856
rect 83100 800 83116 856
rect 83284 800 83392 856
rect 83560 800 83668 856
rect 83836 800 83852 856
rect 84020 800 84128 856
rect 84296 800 84404 856
rect 84572 800 84588 856
rect 84756 800 84864 856
rect 85032 800 85140 856
rect 85308 800 85324 856
rect 85492 800 85600 856
rect 85768 800 85876 856
rect 86044 800 86060 856
rect 86228 800 86336 856
rect 86504 800 86612 856
rect 86780 800 86796 856
rect 86964 800 87072 856
rect 87240 800 87348 856
rect 87516 800 87532 856
rect 87700 800 87808 856
rect 87976 800 88084 856
rect 88252 800 88268 856
rect 88436 800 88544 856
rect 88712 800 88820 856
rect 88988 800 89004 856
rect 89172 800 89280 856
rect 89448 800 89556 856
rect 89724 800 89740 856
rect 89908 800 90016 856
rect 90184 800 90200 856
rect 90368 800 90476 856
rect 90644 800 90752 856
rect 90920 800 90936 856
rect 91104 800 91212 856
rect 91380 800 91488 856
rect 91656 800 91672 856
rect 91840 800 91948 856
rect 92116 800 92224 856
rect 92392 800 92408 856
rect 92576 800 92684 856
rect 92852 800 92960 856
rect 93128 800 93144 856
rect 93312 800 93420 856
rect 93588 800 93696 856
rect 93864 800 93880 856
rect 94048 800 94156 856
rect 94324 800 94432 856
rect 94600 800 94616 856
rect 94784 800 94892 856
rect 95060 800 95168 856
rect 95336 800 95352 856
rect 95520 800 95628 856
rect 95796 800 95904 856
rect 96072 800 96088 856
rect 96256 800 96364 856
rect 96532 800 96640 856
rect 96808 800 96824 856
rect 96992 800 97100 856
rect 97268 800 97376 856
rect 97544 800 97560 856
rect 97728 800 97836 856
rect 98004 800 98112 856
rect 98280 800 98296 856
rect 98464 800 98572 856
rect 98740 800 98848 856
rect 99016 800 99032 856
rect 99200 800 99308 856
rect 99476 800 99584 856
rect 99752 800 99768 856
rect 99936 800 100044 856
rect 100212 800 100320 856
rect 100488 800 100504 856
rect 100672 800 100780 856
rect 100948 800 101056 856
rect 101224 800 101240 856
rect 101408 800 101516 856
rect 101684 800 101792 856
rect 101960 800 101976 856
rect 102144 800 102252 856
rect 102420 800 102528 856
rect 102696 800 102712 856
rect 102880 800 102988 856
rect 103156 800 103264 856
rect 103432 800 103448 856
rect 103616 800 103724 856
rect 103892 800 104000 856
rect 104168 800 104184 856
rect 104352 800 104460 856
rect 104628 800 104736 856
rect 104904 800 104920 856
rect 105088 800 105196 856
rect 105364 800 105380 856
rect 105548 800 105656 856
rect 105824 800 105932 856
rect 106100 800 106116 856
rect 106284 800 106392 856
rect 106560 800 106668 856
rect 106836 800 106852 856
rect 107020 800 107128 856
rect 107296 800 107404 856
rect 107572 800 107588 856
rect 107756 800 107864 856
rect 108032 800 108140 856
rect 108308 800 108324 856
rect 108492 800 108600 856
rect 108768 800 108876 856
rect 109044 800 109060 856
rect 109228 800 109336 856
rect 109504 800 109612 856
rect 109780 800 109796 856
rect 109964 800 110072 856
rect 110240 800 110348 856
rect 110516 800 110532 856
rect 110700 800 110808 856
rect 110976 800 111084 856
rect 111252 800 111268 856
rect 111436 800 111544 856
rect 111712 800 111820 856
rect 111988 800 112004 856
rect 112172 800 112280 856
rect 112448 800 112556 856
rect 112724 800 112740 856
rect 112908 800 113016 856
rect 113184 800 113292 856
rect 113460 800 113476 856
rect 113644 800 113752 856
rect 113920 800 114028 856
rect 114196 800 114212 856
rect 114380 800 114488 856
rect 114656 800 114764 856
rect 114932 800 114948 856
rect 115116 800 115224 856
rect 115392 800 115500 856
rect 115668 800 115684 856
rect 115852 800 115960 856
rect 116128 800 116236 856
rect 116404 800 116420 856
rect 116588 800 116696 856
rect 116864 800 116972 856
rect 117140 800 117156 856
rect 117324 800 117432 856
rect 117600 800 117708 856
rect 117876 800 117892 856
rect 118060 800 118168 856
rect 118336 800 118444 856
rect 118612 800 118628 856
rect 118796 800 118904 856
rect 119072 800 119180 856
rect 119348 800 119364 856
<< obsm3 >>
rect 3679 851 111942 117537
<< metal4 >>
rect 4102 2128 4422 117552
rect 4762 2176 5082 117504
rect 5422 2176 5742 117504
rect 6082 2176 6402 117504
rect 19462 2128 19782 117552
rect 20122 2176 20442 117504
rect 20782 2176 21102 117504
rect 21442 2176 21762 117504
rect 34822 2128 35142 117552
rect 35482 2176 35802 117504
rect 36142 2176 36462 117504
rect 36802 2176 37122 117504
rect 50182 2128 50502 117552
rect 50842 2176 51162 117504
rect 51502 2176 51822 117504
rect 52162 2176 52482 117504
rect 65542 2128 65862 117552
rect 66202 2176 66522 117504
rect 66862 2176 67182 117504
rect 67522 2176 67842 117504
rect 80902 2128 81222 117552
rect 81562 2176 81882 117504
rect 82222 2176 82542 117504
rect 82882 2176 83202 117504
rect 96262 2128 96582 117552
rect 96922 2176 97242 117504
rect 97582 2176 97902 117504
rect 98242 2176 98562 117504
rect 111622 2128 111942 117552
rect 112282 2176 112602 117504
rect 112942 2176 113262 117504
rect 113602 2176 113922 117504
<< obsm4 >>
rect 6577 8331 19382 95165
rect 19862 8331 20042 95165
rect 20522 8331 20702 95165
rect 21182 8331 21362 95165
rect 21842 8331 34742 95165
rect 35222 8331 35402 95165
rect 35882 8331 36062 95165
rect 36542 8331 36722 95165
rect 37202 8331 50102 95165
rect 50582 8331 50762 95165
rect 51242 8331 51422 95165
rect 51902 8331 52082 95165
rect 52562 8331 65462 95165
rect 65942 8331 66122 95165
rect 66602 8331 66782 95165
rect 67262 8331 67442 95165
rect 67922 8331 80427 95165
<< labels >>
rlabel metal2 s 372 119200 428 120000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 31928 119200 31984 120000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 35056 119200 35112 120000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 38184 119200 38240 120000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 41404 119200 41460 120000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 44532 119200 44588 120000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 47660 119200 47716 120000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 50880 119200 50936 120000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 54008 119200 54064 120000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 57136 119200 57192 120000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 60356 119200 60412 120000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 3500 119200 3556 120000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 63484 119200 63540 120000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 66612 119200 66668 120000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 69740 119200 69796 120000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 72960 119200 73016 120000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 76088 119200 76144 120000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 79216 119200 79272 120000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 82436 119200 82492 120000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 85564 119200 85620 120000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 88692 119200 88748 120000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 91912 119200 91968 120000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 6628 119200 6684 120000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 95040 119200 95096 120000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 98168 119200 98224 120000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 101388 119200 101444 120000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 104516 119200 104572 120000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 107644 119200 107700 120000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 110864 119200 110920 120000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 113992 119200 114048 120000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 117120 119200 117176 120000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 9756 119200 9812 120000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 12976 119200 13032 120000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 16104 119200 16160 120000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 19232 119200 19288 120000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 22452 119200 22508 120000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 25580 119200 25636 120000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 28708 119200 28764 120000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1384 119200 1440 120000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 32940 119200 32996 120000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 36068 119200 36124 120000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 39288 119200 39344 120000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 42416 119200 42472 120000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 45544 119200 45600 120000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 48764 119200 48820 120000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 51892 119200 51948 120000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 55020 119200 55076 120000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 58240 119200 58296 120000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 61368 119200 61424 120000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 4512 119200 4568 120000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 64496 119200 64552 120000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 67716 119200 67772 120000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 70844 119200 70900 120000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 73972 119200 74028 120000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 77192 119200 77248 120000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 80320 119200 80376 120000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 83448 119200 83504 120000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 86576 119200 86632 120000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 89796 119200 89852 120000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 92924 119200 92980 120000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 7732 119200 7788 120000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 96052 119200 96108 120000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 99272 119200 99328 120000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 102400 119200 102456 120000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 105528 119200 105584 120000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 108748 119200 108804 120000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 111876 119200 111932 120000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 115004 119200 115060 120000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 118224 119200 118280 120000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 10860 119200 10916 120000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 13988 119200 14044 120000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 17208 119200 17264 120000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 20336 119200 20392 120000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 23464 119200 23520 120000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 26592 119200 26648 120000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 29812 119200 29868 120000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 2396 119200 2452 120000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 34044 119200 34100 120000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 37172 119200 37228 120000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 40300 119200 40356 120000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 43428 119200 43484 120000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 46648 119200 46704 120000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 49776 119200 49832 120000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 52904 119200 52960 120000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 56124 119200 56180 120000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 59252 119200 59308 120000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 62380 119200 62436 120000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 5616 119200 5672 120000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 65600 119200 65656 120000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 68728 119200 68784 120000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 71856 119200 71912 120000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 75076 119200 75132 120000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 78204 119200 78260 120000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 81332 119200 81388 120000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 84552 119200 84608 120000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 87680 119200 87736 120000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 90808 119200 90864 120000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 94028 119200 94084 120000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 8744 119200 8800 120000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 97156 119200 97212 120000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 100284 119200 100340 120000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 103412 119200 103468 120000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 106632 119200 106688 120000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 109760 119200 109816 120000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 112888 119200 112944 120000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 116108 119200 116164 120000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 119236 119200 119292 120000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 11872 119200 11928 120000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 15092 119200 15148 120000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 18220 119200 18276 120000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 21348 119200 21404 120000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 24568 119200 24624 120000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 27696 119200 27752 120000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 30824 119200 30880 120000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 25948 0 26004 800 6 la_data_in[0]
port 115 nsew signal input
rlabel metal2 s 99364 0 99420 800 6 la_data_in[100]
port 116 nsew signal input
rlabel metal2 s 100100 0 100156 800 6 la_data_in[101]
port 117 nsew signal input
rlabel metal2 s 100836 0 100892 800 6 la_data_in[102]
port 118 nsew signal input
rlabel metal2 s 101572 0 101628 800 6 la_data_in[103]
port 119 nsew signal input
rlabel metal2 s 102308 0 102364 800 6 la_data_in[104]
port 120 nsew signal input
rlabel metal2 s 103044 0 103100 800 6 la_data_in[105]
port 121 nsew signal input
rlabel metal2 s 103780 0 103836 800 6 la_data_in[106]
port 122 nsew signal input
rlabel metal2 s 104516 0 104572 800 6 la_data_in[107]
port 123 nsew signal input
rlabel metal2 s 105252 0 105308 800 6 la_data_in[108]
port 124 nsew signal input
rlabel metal2 s 105988 0 106044 800 6 la_data_in[109]
port 125 nsew signal input
rlabel metal2 s 33216 0 33272 800 6 la_data_in[10]
port 126 nsew signal input
rlabel metal2 s 106724 0 106780 800 6 la_data_in[110]
port 127 nsew signal input
rlabel metal2 s 107460 0 107516 800 6 la_data_in[111]
port 128 nsew signal input
rlabel metal2 s 108196 0 108252 800 6 la_data_in[112]
port 129 nsew signal input
rlabel metal2 s 108932 0 108988 800 6 la_data_in[113]
port 130 nsew signal input
rlabel metal2 s 109668 0 109724 800 6 la_data_in[114]
port 131 nsew signal input
rlabel metal2 s 110404 0 110460 800 6 la_data_in[115]
port 132 nsew signal input
rlabel metal2 s 111140 0 111196 800 6 la_data_in[116]
port 133 nsew signal input
rlabel metal2 s 111876 0 111932 800 6 la_data_in[117]
port 134 nsew signal input
rlabel metal2 s 112612 0 112668 800 6 la_data_in[118]
port 135 nsew signal input
rlabel metal2 s 113348 0 113404 800 6 la_data_in[119]
port 136 nsew signal input
rlabel metal2 s 33952 0 34008 800 6 la_data_in[11]
port 137 nsew signal input
rlabel metal2 s 114084 0 114140 800 6 la_data_in[120]
port 138 nsew signal input
rlabel metal2 s 114820 0 114876 800 6 la_data_in[121]
port 139 nsew signal input
rlabel metal2 s 115556 0 115612 800 6 la_data_in[122]
port 140 nsew signal input
rlabel metal2 s 116292 0 116348 800 6 la_data_in[123]
port 141 nsew signal input
rlabel metal2 s 117028 0 117084 800 6 la_data_in[124]
port 142 nsew signal input
rlabel metal2 s 117764 0 117820 800 6 la_data_in[125]
port 143 nsew signal input
rlabel metal2 s 118500 0 118556 800 6 la_data_in[126]
port 144 nsew signal input
rlabel metal2 s 119236 0 119292 800 6 la_data_in[127]
port 145 nsew signal input
rlabel metal2 s 34688 0 34744 800 6 la_data_in[12]
port 146 nsew signal input
rlabel metal2 s 35424 0 35480 800 6 la_data_in[13]
port 147 nsew signal input
rlabel metal2 s 36160 0 36216 800 6 la_data_in[14]
port 148 nsew signal input
rlabel metal2 s 36896 0 36952 800 6 la_data_in[15]
port 149 nsew signal input
rlabel metal2 s 37632 0 37688 800 6 la_data_in[16]
port 150 nsew signal input
rlabel metal2 s 38368 0 38424 800 6 la_data_in[17]
port 151 nsew signal input
rlabel metal2 s 39104 0 39160 800 6 la_data_in[18]
port 152 nsew signal input
rlabel metal2 s 39840 0 39896 800 6 la_data_in[19]
port 153 nsew signal input
rlabel metal2 s 26684 0 26740 800 6 la_data_in[1]
port 154 nsew signal input
rlabel metal2 s 40576 0 40632 800 6 la_data_in[20]
port 155 nsew signal input
rlabel metal2 s 41312 0 41368 800 6 la_data_in[21]
port 156 nsew signal input
rlabel metal2 s 42048 0 42104 800 6 la_data_in[22]
port 157 nsew signal input
rlabel metal2 s 42784 0 42840 800 6 la_data_in[23]
port 158 nsew signal input
rlabel metal2 s 43520 0 43576 800 6 la_data_in[24]
port 159 nsew signal input
rlabel metal2 s 44256 0 44312 800 6 la_data_in[25]
port 160 nsew signal input
rlabel metal2 s 44992 0 45048 800 6 la_data_in[26]
port 161 nsew signal input
rlabel metal2 s 45728 0 45784 800 6 la_data_in[27]
port 162 nsew signal input
rlabel metal2 s 46464 0 46520 800 6 la_data_in[28]
port 163 nsew signal input
rlabel metal2 s 47200 0 47256 800 6 la_data_in[29]
port 164 nsew signal input
rlabel metal2 s 27420 0 27476 800 6 la_data_in[2]
port 165 nsew signal input
rlabel metal2 s 47936 0 47992 800 6 la_data_in[30]
port 166 nsew signal input
rlabel metal2 s 48672 0 48728 800 6 la_data_in[31]
port 167 nsew signal input
rlabel metal2 s 49408 0 49464 800 6 la_data_in[32]
port 168 nsew signal input
rlabel metal2 s 50144 0 50200 800 6 la_data_in[33]
port 169 nsew signal input
rlabel metal2 s 50880 0 50936 800 6 la_data_in[34]
port 170 nsew signal input
rlabel metal2 s 51616 0 51672 800 6 la_data_in[35]
port 171 nsew signal input
rlabel metal2 s 52352 0 52408 800 6 la_data_in[36]
port 172 nsew signal input
rlabel metal2 s 53088 0 53144 800 6 la_data_in[37]
port 173 nsew signal input
rlabel metal2 s 53824 0 53880 800 6 la_data_in[38]
port 174 nsew signal input
rlabel metal2 s 54560 0 54616 800 6 la_data_in[39]
port 175 nsew signal input
rlabel metal2 s 28156 0 28212 800 6 la_data_in[3]
port 176 nsew signal input
rlabel metal2 s 55296 0 55352 800 6 la_data_in[40]
port 177 nsew signal input
rlabel metal2 s 56032 0 56088 800 6 la_data_in[41]
port 178 nsew signal input
rlabel metal2 s 56768 0 56824 800 6 la_data_in[42]
port 179 nsew signal input
rlabel metal2 s 57504 0 57560 800 6 la_data_in[43]
port 180 nsew signal input
rlabel metal2 s 58240 0 58296 800 6 la_data_in[44]
port 181 nsew signal input
rlabel metal2 s 58976 0 59032 800 6 la_data_in[45]
port 182 nsew signal input
rlabel metal2 s 59712 0 59768 800 6 la_data_in[46]
port 183 nsew signal input
rlabel metal2 s 60448 0 60504 800 6 la_data_in[47]
port 184 nsew signal input
rlabel metal2 s 61184 0 61240 800 6 la_data_in[48]
port 185 nsew signal input
rlabel metal2 s 61920 0 61976 800 6 la_data_in[49]
port 186 nsew signal input
rlabel metal2 s 28892 0 28948 800 6 la_data_in[4]
port 187 nsew signal input
rlabel metal2 s 62656 0 62712 800 6 la_data_in[50]
port 188 nsew signal input
rlabel metal2 s 63392 0 63448 800 6 la_data_in[51]
port 189 nsew signal input
rlabel metal2 s 64128 0 64184 800 6 la_data_in[52]
port 190 nsew signal input
rlabel metal2 s 64864 0 64920 800 6 la_data_in[53]
port 191 nsew signal input
rlabel metal2 s 65600 0 65656 800 6 la_data_in[54]
port 192 nsew signal input
rlabel metal2 s 66336 0 66392 800 6 la_data_in[55]
port 193 nsew signal input
rlabel metal2 s 67072 0 67128 800 6 la_data_in[56]
port 194 nsew signal input
rlabel metal2 s 67808 0 67864 800 6 la_data_in[57]
port 195 nsew signal input
rlabel metal2 s 68544 0 68600 800 6 la_data_in[58]
port 196 nsew signal input
rlabel metal2 s 69280 0 69336 800 6 la_data_in[59]
port 197 nsew signal input
rlabel metal2 s 29628 0 29684 800 6 la_data_in[5]
port 198 nsew signal input
rlabel metal2 s 70016 0 70072 800 6 la_data_in[60]
port 199 nsew signal input
rlabel metal2 s 70752 0 70808 800 6 la_data_in[61]
port 200 nsew signal input
rlabel metal2 s 71488 0 71544 800 6 la_data_in[62]
port 201 nsew signal input
rlabel metal2 s 72224 0 72280 800 6 la_data_in[63]
port 202 nsew signal input
rlabel metal2 s 72960 0 73016 800 6 la_data_in[64]
port 203 nsew signal input
rlabel metal2 s 73696 0 73752 800 6 la_data_in[65]
port 204 nsew signal input
rlabel metal2 s 74432 0 74488 800 6 la_data_in[66]
port 205 nsew signal input
rlabel metal2 s 75076 0 75132 800 6 la_data_in[67]
port 206 nsew signal input
rlabel metal2 s 75812 0 75868 800 6 la_data_in[68]
port 207 nsew signal input
rlabel metal2 s 76548 0 76604 800 6 la_data_in[69]
port 208 nsew signal input
rlabel metal2 s 30272 0 30328 800 6 la_data_in[6]
port 209 nsew signal input
rlabel metal2 s 77284 0 77340 800 6 la_data_in[70]
port 210 nsew signal input
rlabel metal2 s 78020 0 78076 800 6 la_data_in[71]
port 211 nsew signal input
rlabel metal2 s 78756 0 78812 800 6 la_data_in[72]
port 212 nsew signal input
rlabel metal2 s 79492 0 79548 800 6 la_data_in[73]
port 213 nsew signal input
rlabel metal2 s 80228 0 80284 800 6 la_data_in[74]
port 214 nsew signal input
rlabel metal2 s 80964 0 81020 800 6 la_data_in[75]
port 215 nsew signal input
rlabel metal2 s 81700 0 81756 800 6 la_data_in[76]
port 216 nsew signal input
rlabel metal2 s 82436 0 82492 800 6 la_data_in[77]
port 217 nsew signal input
rlabel metal2 s 83172 0 83228 800 6 la_data_in[78]
port 218 nsew signal input
rlabel metal2 s 83908 0 83964 800 6 la_data_in[79]
port 219 nsew signal input
rlabel metal2 s 31008 0 31064 800 6 la_data_in[7]
port 220 nsew signal input
rlabel metal2 s 84644 0 84700 800 6 la_data_in[80]
port 221 nsew signal input
rlabel metal2 s 85380 0 85436 800 6 la_data_in[81]
port 222 nsew signal input
rlabel metal2 s 86116 0 86172 800 6 la_data_in[82]
port 223 nsew signal input
rlabel metal2 s 86852 0 86908 800 6 la_data_in[83]
port 224 nsew signal input
rlabel metal2 s 87588 0 87644 800 6 la_data_in[84]
port 225 nsew signal input
rlabel metal2 s 88324 0 88380 800 6 la_data_in[85]
port 226 nsew signal input
rlabel metal2 s 89060 0 89116 800 6 la_data_in[86]
port 227 nsew signal input
rlabel metal2 s 89796 0 89852 800 6 la_data_in[87]
port 228 nsew signal input
rlabel metal2 s 90532 0 90588 800 6 la_data_in[88]
port 229 nsew signal input
rlabel metal2 s 91268 0 91324 800 6 la_data_in[89]
port 230 nsew signal input
rlabel metal2 s 31744 0 31800 800 6 la_data_in[8]
port 231 nsew signal input
rlabel metal2 s 92004 0 92060 800 6 la_data_in[90]
port 232 nsew signal input
rlabel metal2 s 92740 0 92796 800 6 la_data_in[91]
port 233 nsew signal input
rlabel metal2 s 93476 0 93532 800 6 la_data_in[92]
port 234 nsew signal input
rlabel metal2 s 94212 0 94268 800 6 la_data_in[93]
port 235 nsew signal input
rlabel metal2 s 94948 0 95004 800 6 la_data_in[94]
port 236 nsew signal input
rlabel metal2 s 95684 0 95740 800 6 la_data_in[95]
port 237 nsew signal input
rlabel metal2 s 96420 0 96476 800 6 la_data_in[96]
port 238 nsew signal input
rlabel metal2 s 97156 0 97212 800 6 la_data_in[97]
port 239 nsew signal input
rlabel metal2 s 97892 0 97948 800 6 la_data_in[98]
port 240 nsew signal input
rlabel metal2 s 98628 0 98684 800 6 la_data_in[99]
port 241 nsew signal input
rlabel metal2 s 32480 0 32536 800 6 la_data_in[9]
port 242 nsew signal input
rlabel metal2 s 26132 0 26188 800 6 la_data_out[0]
port 243 nsew signal output
rlabel metal2 s 99640 0 99696 800 6 la_data_out[100]
port 244 nsew signal output
rlabel metal2 s 100376 0 100432 800 6 la_data_out[101]
port 245 nsew signal output
rlabel metal2 s 101112 0 101168 800 6 la_data_out[102]
port 246 nsew signal output
rlabel metal2 s 101848 0 101904 800 6 la_data_out[103]
port 247 nsew signal output
rlabel metal2 s 102584 0 102640 800 6 la_data_out[104]
port 248 nsew signal output
rlabel metal2 s 103320 0 103376 800 6 la_data_out[105]
port 249 nsew signal output
rlabel metal2 s 104056 0 104112 800 6 la_data_out[106]
port 250 nsew signal output
rlabel metal2 s 104792 0 104848 800 6 la_data_out[107]
port 251 nsew signal output
rlabel metal2 s 105436 0 105492 800 6 la_data_out[108]
port 252 nsew signal output
rlabel metal2 s 106172 0 106228 800 6 la_data_out[109]
port 253 nsew signal output
rlabel metal2 s 33492 0 33548 800 6 la_data_out[10]
port 254 nsew signal output
rlabel metal2 s 106908 0 106964 800 6 la_data_out[110]
port 255 nsew signal output
rlabel metal2 s 107644 0 107700 800 6 la_data_out[111]
port 256 nsew signal output
rlabel metal2 s 108380 0 108436 800 6 la_data_out[112]
port 257 nsew signal output
rlabel metal2 s 109116 0 109172 800 6 la_data_out[113]
port 258 nsew signal output
rlabel metal2 s 109852 0 109908 800 6 la_data_out[114]
port 259 nsew signal output
rlabel metal2 s 110588 0 110644 800 6 la_data_out[115]
port 260 nsew signal output
rlabel metal2 s 111324 0 111380 800 6 la_data_out[116]
port 261 nsew signal output
rlabel metal2 s 112060 0 112116 800 6 la_data_out[117]
port 262 nsew signal output
rlabel metal2 s 112796 0 112852 800 6 la_data_out[118]
port 263 nsew signal output
rlabel metal2 s 113532 0 113588 800 6 la_data_out[119]
port 264 nsew signal output
rlabel metal2 s 34228 0 34284 800 6 la_data_out[11]
port 265 nsew signal output
rlabel metal2 s 114268 0 114324 800 6 la_data_out[120]
port 266 nsew signal output
rlabel metal2 s 115004 0 115060 800 6 la_data_out[121]
port 267 nsew signal output
rlabel metal2 s 115740 0 115796 800 6 la_data_out[122]
port 268 nsew signal output
rlabel metal2 s 116476 0 116532 800 6 la_data_out[123]
port 269 nsew signal output
rlabel metal2 s 117212 0 117268 800 6 la_data_out[124]
port 270 nsew signal output
rlabel metal2 s 117948 0 118004 800 6 la_data_out[125]
port 271 nsew signal output
rlabel metal2 s 118684 0 118740 800 6 la_data_out[126]
port 272 nsew signal output
rlabel metal2 s 119420 0 119476 800 6 la_data_out[127]
port 273 nsew signal output
rlabel metal2 s 34964 0 35020 800 6 la_data_out[12]
port 274 nsew signal output
rlabel metal2 s 35700 0 35756 800 6 la_data_out[13]
port 275 nsew signal output
rlabel metal2 s 36436 0 36492 800 6 la_data_out[14]
port 276 nsew signal output
rlabel metal2 s 37172 0 37228 800 6 la_data_out[15]
port 277 nsew signal output
rlabel metal2 s 37908 0 37964 800 6 la_data_out[16]
port 278 nsew signal output
rlabel metal2 s 38644 0 38700 800 6 la_data_out[17]
port 279 nsew signal output
rlabel metal2 s 39380 0 39436 800 6 la_data_out[18]
port 280 nsew signal output
rlabel metal2 s 40116 0 40172 800 6 la_data_out[19]
port 281 nsew signal output
rlabel metal2 s 26868 0 26924 800 6 la_data_out[1]
port 282 nsew signal output
rlabel metal2 s 40852 0 40908 800 6 la_data_out[20]
port 283 nsew signal output
rlabel metal2 s 41588 0 41644 800 6 la_data_out[21]
port 284 nsew signal output
rlabel metal2 s 42324 0 42380 800 6 la_data_out[22]
port 285 nsew signal output
rlabel metal2 s 43060 0 43116 800 6 la_data_out[23]
port 286 nsew signal output
rlabel metal2 s 43796 0 43852 800 6 la_data_out[24]
port 287 nsew signal output
rlabel metal2 s 44532 0 44588 800 6 la_data_out[25]
port 288 nsew signal output
rlabel metal2 s 45268 0 45324 800 6 la_data_out[26]
port 289 nsew signal output
rlabel metal2 s 46004 0 46060 800 6 la_data_out[27]
port 290 nsew signal output
rlabel metal2 s 46740 0 46796 800 6 la_data_out[28]
port 291 nsew signal output
rlabel metal2 s 47476 0 47532 800 6 la_data_out[29]
port 292 nsew signal output
rlabel metal2 s 27604 0 27660 800 6 la_data_out[2]
port 293 nsew signal output
rlabel metal2 s 48212 0 48268 800 6 la_data_out[30]
port 294 nsew signal output
rlabel metal2 s 48948 0 49004 800 6 la_data_out[31]
port 295 nsew signal output
rlabel metal2 s 49684 0 49740 800 6 la_data_out[32]
port 296 nsew signal output
rlabel metal2 s 50420 0 50476 800 6 la_data_out[33]
port 297 nsew signal output
rlabel metal2 s 51156 0 51212 800 6 la_data_out[34]
port 298 nsew signal output
rlabel metal2 s 51892 0 51948 800 6 la_data_out[35]
port 299 nsew signal output
rlabel metal2 s 52628 0 52684 800 6 la_data_out[36]
port 300 nsew signal output
rlabel metal2 s 53364 0 53420 800 6 la_data_out[37]
port 301 nsew signal output
rlabel metal2 s 54100 0 54156 800 6 la_data_out[38]
port 302 nsew signal output
rlabel metal2 s 54836 0 54892 800 6 la_data_out[39]
port 303 nsew signal output
rlabel metal2 s 28340 0 28396 800 6 la_data_out[3]
port 304 nsew signal output
rlabel metal2 s 55572 0 55628 800 6 la_data_out[40]
port 305 nsew signal output
rlabel metal2 s 56308 0 56364 800 6 la_data_out[41]
port 306 nsew signal output
rlabel metal2 s 57044 0 57100 800 6 la_data_out[42]
port 307 nsew signal output
rlabel metal2 s 57780 0 57836 800 6 la_data_out[43]
port 308 nsew signal output
rlabel metal2 s 58516 0 58572 800 6 la_data_out[44]
port 309 nsew signal output
rlabel metal2 s 59252 0 59308 800 6 la_data_out[45]
port 310 nsew signal output
rlabel metal2 s 59988 0 60044 800 6 la_data_out[46]
port 311 nsew signal output
rlabel metal2 s 60632 0 60688 800 6 la_data_out[47]
port 312 nsew signal output
rlabel metal2 s 61368 0 61424 800 6 la_data_out[48]
port 313 nsew signal output
rlabel metal2 s 62104 0 62160 800 6 la_data_out[49]
port 314 nsew signal output
rlabel metal2 s 29076 0 29132 800 6 la_data_out[4]
port 315 nsew signal output
rlabel metal2 s 62840 0 62896 800 6 la_data_out[50]
port 316 nsew signal output
rlabel metal2 s 63576 0 63632 800 6 la_data_out[51]
port 317 nsew signal output
rlabel metal2 s 64312 0 64368 800 6 la_data_out[52]
port 318 nsew signal output
rlabel metal2 s 65048 0 65104 800 6 la_data_out[53]
port 319 nsew signal output
rlabel metal2 s 65784 0 65840 800 6 la_data_out[54]
port 320 nsew signal output
rlabel metal2 s 66520 0 66576 800 6 la_data_out[55]
port 321 nsew signal output
rlabel metal2 s 67256 0 67312 800 6 la_data_out[56]
port 322 nsew signal output
rlabel metal2 s 67992 0 68048 800 6 la_data_out[57]
port 323 nsew signal output
rlabel metal2 s 68728 0 68784 800 6 la_data_out[58]
port 324 nsew signal output
rlabel metal2 s 69464 0 69520 800 6 la_data_out[59]
port 325 nsew signal output
rlabel metal2 s 29812 0 29868 800 6 la_data_out[5]
port 326 nsew signal output
rlabel metal2 s 70200 0 70256 800 6 la_data_out[60]
port 327 nsew signal output
rlabel metal2 s 70936 0 70992 800 6 la_data_out[61]
port 328 nsew signal output
rlabel metal2 s 71672 0 71728 800 6 la_data_out[62]
port 329 nsew signal output
rlabel metal2 s 72408 0 72464 800 6 la_data_out[63]
port 330 nsew signal output
rlabel metal2 s 73144 0 73200 800 6 la_data_out[64]
port 331 nsew signal output
rlabel metal2 s 73880 0 73936 800 6 la_data_out[65]
port 332 nsew signal output
rlabel metal2 s 74616 0 74672 800 6 la_data_out[66]
port 333 nsew signal output
rlabel metal2 s 75352 0 75408 800 6 la_data_out[67]
port 334 nsew signal output
rlabel metal2 s 76088 0 76144 800 6 la_data_out[68]
port 335 nsew signal output
rlabel metal2 s 76824 0 76880 800 6 la_data_out[69]
port 336 nsew signal output
rlabel metal2 s 30548 0 30604 800 6 la_data_out[6]
port 337 nsew signal output
rlabel metal2 s 77560 0 77616 800 6 la_data_out[70]
port 338 nsew signal output
rlabel metal2 s 78296 0 78352 800 6 la_data_out[71]
port 339 nsew signal output
rlabel metal2 s 79032 0 79088 800 6 la_data_out[72]
port 340 nsew signal output
rlabel metal2 s 79768 0 79824 800 6 la_data_out[73]
port 341 nsew signal output
rlabel metal2 s 80504 0 80560 800 6 la_data_out[74]
port 342 nsew signal output
rlabel metal2 s 81240 0 81296 800 6 la_data_out[75]
port 343 nsew signal output
rlabel metal2 s 81976 0 82032 800 6 la_data_out[76]
port 344 nsew signal output
rlabel metal2 s 82712 0 82768 800 6 la_data_out[77]
port 345 nsew signal output
rlabel metal2 s 83448 0 83504 800 6 la_data_out[78]
port 346 nsew signal output
rlabel metal2 s 84184 0 84240 800 6 la_data_out[79]
port 347 nsew signal output
rlabel metal2 s 31284 0 31340 800 6 la_data_out[7]
port 348 nsew signal output
rlabel metal2 s 84920 0 84976 800 6 la_data_out[80]
port 349 nsew signal output
rlabel metal2 s 85656 0 85712 800 6 la_data_out[81]
port 350 nsew signal output
rlabel metal2 s 86392 0 86448 800 6 la_data_out[82]
port 351 nsew signal output
rlabel metal2 s 87128 0 87184 800 6 la_data_out[83]
port 352 nsew signal output
rlabel metal2 s 87864 0 87920 800 6 la_data_out[84]
port 353 nsew signal output
rlabel metal2 s 88600 0 88656 800 6 la_data_out[85]
port 354 nsew signal output
rlabel metal2 s 89336 0 89392 800 6 la_data_out[86]
port 355 nsew signal output
rlabel metal2 s 90072 0 90128 800 6 la_data_out[87]
port 356 nsew signal output
rlabel metal2 s 90808 0 90864 800 6 la_data_out[88]
port 357 nsew signal output
rlabel metal2 s 91544 0 91600 800 6 la_data_out[89]
port 358 nsew signal output
rlabel metal2 s 32020 0 32076 800 6 la_data_out[8]
port 359 nsew signal output
rlabel metal2 s 92280 0 92336 800 6 la_data_out[90]
port 360 nsew signal output
rlabel metal2 s 93016 0 93072 800 6 la_data_out[91]
port 361 nsew signal output
rlabel metal2 s 93752 0 93808 800 6 la_data_out[92]
port 362 nsew signal output
rlabel metal2 s 94488 0 94544 800 6 la_data_out[93]
port 363 nsew signal output
rlabel metal2 s 95224 0 95280 800 6 la_data_out[94]
port 364 nsew signal output
rlabel metal2 s 95960 0 96016 800 6 la_data_out[95]
port 365 nsew signal output
rlabel metal2 s 96696 0 96752 800 6 la_data_out[96]
port 366 nsew signal output
rlabel metal2 s 97432 0 97488 800 6 la_data_out[97]
port 367 nsew signal output
rlabel metal2 s 98168 0 98224 800 6 la_data_out[98]
port 368 nsew signal output
rlabel metal2 s 98904 0 98960 800 6 la_data_out[99]
port 369 nsew signal output
rlabel metal2 s 32756 0 32812 800 6 la_data_out[9]
port 370 nsew signal output
rlabel metal2 s 26408 0 26464 800 6 la_oen[0]
port 371 nsew signal input
rlabel metal2 s 99824 0 99880 800 6 la_oen[100]
port 372 nsew signal input
rlabel metal2 s 100560 0 100616 800 6 la_oen[101]
port 373 nsew signal input
rlabel metal2 s 101296 0 101352 800 6 la_oen[102]
port 374 nsew signal input
rlabel metal2 s 102032 0 102088 800 6 la_oen[103]
port 375 nsew signal input
rlabel metal2 s 102768 0 102824 800 6 la_oen[104]
port 376 nsew signal input
rlabel metal2 s 103504 0 103560 800 6 la_oen[105]
port 377 nsew signal input
rlabel metal2 s 104240 0 104296 800 6 la_oen[106]
port 378 nsew signal input
rlabel metal2 s 104976 0 105032 800 6 la_oen[107]
port 379 nsew signal input
rlabel metal2 s 105712 0 105768 800 6 la_oen[108]
port 380 nsew signal input
rlabel metal2 s 106448 0 106504 800 6 la_oen[109]
port 381 nsew signal input
rlabel metal2 s 33768 0 33824 800 6 la_oen[10]
port 382 nsew signal input
rlabel metal2 s 107184 0 107240 800 6 la_oen[110]
port 383 nsew signal input
rlabel metal2 s 107920 0 107976 800 6 la_oen[111]
port 384 nsew signal input
rlabel metal2 s 108656 0 108712 800 6 la_oen[112]
port 385 nsew signal input
rlabel metal2 s 109392 0 109448 800 6 la_oen[113]
port 386 nsew signal input
rlabel metal2 s 110128 0 110184 800 6 la_oen[114]
port 387 nsew signal input
rlabel metal2 s 110864 0 110920 800 6 la_oen[115]
port 388 nsew signal input
rlabel metal2 s 111600 0 111656 800 6 la_oen[116]
port 389 nsew signal input
rlabel metal2 s 112336 0 112392 800 6 la_oen[117]
port 390 nsew signal input
rlabel metal2 s 113072 0 113128 800 6 la_oen[118]
port 391 nsew signal input
rlabel metal2 s 113808 0 113864 800 6 la_oen[119]
port 392 nsew signal input
rlabel metal2 s 34504 0 34560 800 6 la_oen[11]
port 393 nsew signal input
rlabel metal2 s 114544 0 114600 800 6 la_oen[120]
port 394 nsew signal input
rlabel metal2 s 115280 0 115336 800 6 la_oen[121]
port 395 nsew signal input
rlabel metal2 s 116016 0 116072 800 6 la_oen[122]
port 396 nsew signal input
rlabel metal2 s 116752 0 116808 800 6 la_oen[123]
port 397 nsew signal input
rlabel metal2 s 117488 0 117544 800 6 la_oen[124]
port 398 nsew signal input
rlabel metal2 s 118224 0 118280 800 6 la_oen[125]
port 399 nsew signal input
rlabel metal2 s 118960 0 119016 800 6 la_oen[126]
port 400 nsew signal input
rlabel metal2 s 119696 0 119752 800 6 la_oen[127]
port 401 nsew signal input
rlabel metal2 s 35240 0 35296 800 6 la_oen[12]
port 402 nsew signal input
rlabel metal2 s 35976 0 36032 800 6 la_oen[13]
port 403 nsew signal input
rlabel metal2 s 36712 0 36768 800 6 la_oen[14]
port 404 nsew signal input
rlabel metal2 s 37448 0 37504 800 6 la_oen[15]
port 405 nsew signal input
rlabel metal2 s 38184 0 38240 800 6 la_oen[16]
port 406 nsew signal input
rlabel metal2 s 38920 0 38976 800 6 la_oen[17]
port 407 nsew signal input
rlabel metal2 s 39656 0 39712 800 6 la_oen[18]
port 408 nsew signal input
rlabel metal2 s 40392 0 40448 800 6 la_oen[19]
port 409 nsew signal input
rlabel metal2 s 27144 0 27200 800 6 la_oen[1]
port 410 nsew signal input
rlabel metal2 s 41128 0 41184 800 6 la_oen[20]
port 411 nsew signal input
rlabel metal2 s 41864 0 41920 800 6 la_oen[21]
port 412 nsew signal input
rlabel metal2 s 42600 0 42656 800 6 la_oen[22]
port 413 nsew signal input
rlabel metal2 s 43336 0 43392 800 6 la_oen[23]
port 414 nsew signal input
rlabel metal2 s 44072 0 44128 800 6 la_oen[24]
port 415 nsew signal input
rlabel metal2 s 44808 0 44864 800 6 la_oen[25]
port 416 nsew signal input
rlabel metal2 s 45452 0 45508 800 6 la_oen[26]
port 417 nsew signal input
rlabel metal2 s 46188 0 46244 800 6 la_oen[27]
port 418 nsew signal input
rlabel metal2 s 46924 0 46980 800 6 la_oen[28]
port 419 nsew signal input
rlabel metal2 s 47660 0 47716 800 6 la_oen[29]
port 420 nsew signal input
rlabel metal2 s 27880 0 27936 800 6 la_oen[2]
port 421 nsew signal input
rlabel metal2 s 48396 0 48452 800 6 la_oen[30]
port 422 nsew signal input
rlabel metal2 s 49132 0 49188 800 6 la_oen[31]
port 423 nsew signal input
rlabel metal2 s 49868 0 49924 800 6 la_oen[32]
port 424 nsew signal input
rlabel metal2 s 50604 0 50660 800 6 la_oen[33]
port 425 nsew signal input
rlabel metal2 s 51340 0 51396 800 6 la_oen[34]
port 426 nsew signal input
rlabel metal2 s 52076 0 52132 800 6 la_oen[35]
port 427 nsew signal input
rlabel metal2 s 52812 0 52868 800 6 la_oen[36]
port 428 nsew signal input
rlabel metal2 s 53548 0 53604 800 6 la_oen[37]
port 429 nsew signal input
rlabel metal2 s 54284 0 54340 800 6 la_oen[38]
port 430 nsew signal input
rlabel metal2 s 55020 0 55076 800 6 la_oen[39]
port 431 nsew signal input
rlabel metal2 s 28616 0 28672 800 6 la_oen[3]
port 432 nsew signal input
rlabel metal2 s 55756 0 55812 800 6 la_oen[40]
port 433 nsew signal input
rlabel metal2 s 56492 0 56548 800 6 la_oen[41]
port 434 nsew signal input
rlabel metal2 s 57228 0 57284 800 6 la_oen[42]
port 435 nsew signal input
rlabel metal2 s 57964 0 58020 800 6 la_oen[43]
port 436 nsew signal input
rlabel metal2 s 58700 0 58756 800 6 la_oen[44]
port 437 nsew signal input
rlabel metal2 s 59436 0 59492 800 6 la_oen[45]
port 438 nsew signal input
rlabel metal2 s 60172 0 60228 800 6 la_oen[46]
port 439 nsew signal input
rlabel metal2 s 60908 0 60964 800 6 la_oen[47]
port 440 nsew signal input
rlabel metal2 s 61644 0 61700 800 6 la_oen[48]
port 441 nsew signal input
rlabel metal2 s 62380 0 62436 800 6 la_oen[49]
port 442 nsew signal input
rlabel metal2 s 29352 0 29408 800 6 la_oen[4]
port 443 nsew signal input
rlabel metal2 s 63116 0 63172 800 6 la_oen[50]
port 444 nsew signal input
rlabel metal2 s 63852 0 63908 800 6 la_oen[51]
port 445 nsew signal input
rlabel metal2 s 64588 0 64644 800 6 la_oen[52]
port 446 nsew signal input
rlabel metal2 s 65324 0 65380 800 6 la_oen[53]
port 447 nsew signal input
rlabel metal2 s 66060 0 66116 800 6 la_oen[54]
port 448 nsew signal input
rlabel metal2 s 66796 0 66852 800 6 la_oen[55]
port 449 nsew signal input
rlabel metal2 s 67532 0 67588 800 6 la_oen[56]
port 450 nsew signal input
rlabel metal2 s 68268 0 68324 800 6 la_oen[57]
port 451 nsew signal input
rlabel metal2 s 69004 0 69060 800 6 la_oen[58]
port 452 nsew signal input
rlabel metal2 s 69740 0 69796 800 6 la_oen[59]
port 453 nsew signal input
rlabel metal2 s 30088 0 30144 800 6 la_oen[5]
port 454 nsew signal input
rlabel metal2 s 70476 0 70532 800 6 la_oen[60]
port 455 nsew signal input
rlabel metal2 s 71212 0 71268 800 6 la_oen[61]
port 456 nsew signal input
rlabel metal2 s 71948 0 72004 800 6 la_oen[62]
port 457 nsew signal input
rlabel metal2 s 72684 0 72740 800 6 la_oen[63]
port 458 nsew signal input
rlabel metal2 s 73420 0 73476 800 6 la_oen[64]
port 459 nsew signal input
rlabel metal2 s 74156 0 74212 800 6 la_oen[65]
port 460 nsew signal input
rlabel metal2 s 74892 0 74948 800 6 la_oen[66]
port 461 nsew signal input
rlabel metal2 s 75628 0 75684 800 6 la_oen[67]
port 462 nsew signal input
rlabel metal2 s 76364 0 76420 800 6 la_oen[68]
port 463 nsew signal input
rlabel metal2 s 77100 0 77156 800 6 la_oen[69]
port 464 nsew signal input
rlabel metal2 s 30824 0 30880 800 6 la_oen[6]
port 465 nsew signal input
rlabel metal2 s 77836 0 77892 800 6 la_oen[70]
port 466 nsew signal input
rlabel metal2 s 78572 0 78628 800 6 la_oen[71]
port 467 nsew signal input
rlabel metal2 s 79308 0 79364 800 6 la_oen[72]
port 468 nsew signal input
rlabel metal2 s 80044 0 80100 800 6 la_oen[73]
port 469 nsew signal input
rlabel metal2 s 80780 0 80836 800 6 la_oen[74]
port 470 nsew signal input
rlabel metal2 s 81516 0 81572 800 6 la_oen[75]
port 471 nsew signal input
rlabel metal2 s 82252 0 82308 800 6 la_oen[76]
port 472 nsew signal input
rlabel metal2 s 82988 0 83044 800 6 la_oen[77]
port 473 nsew signal input
rlabel metal2 s 83724 0 83780 800 6 la_oen[78]
port 474 nsew signal input
rlabel metal2 s 84460 0 84516 800 6 la_oen[79]
port 475 nsew signal input
rlabel metal2 s 31560 0 31616 800 6 la_oen[7]
port 476 nsew signal input
rlabel metal2 s 85196 0 85252 800 6 la_oen[80]
port 477 nsew signal input
rlabel metal2 s 85932 0 85988 800 6 la_oen[81]
port 478 nsew signal input
rlabel metal2 s 86668 0 86724 800 6 la_oen[82]
port 479 nsew signal input
rlabel metal2 s 87404 0 87460 800 6 la_oen[83]
port 480 nsew signal input
rlabel metal2 s 88140 0 88196 800 6 la_oen[84]
port 481 nsew signal input
rlabel metal2 s 88876 0 88932 800 6 la_oen[85]
port 482 nsew signal input
rlabel metal2 s 89612 0 89668 800 6 la_oen[86]
port 483 nsew signal input
rlabel metal2 s 90256 0 90312 800 6 la_oen[87]
port 484 nsew signal input
rlabel metal2 s 90992 0 91048 800 6 la_oen[88]
port 485 nsew signal input
rlabel metal2 s 91728 0 91784 800 6 la_oen[89]
port 486 nsew signal input
rlabel metal2 s 32296 0 32352 800 6 la_oen[8]
port 487 nsew signal input
rlabel metal2 s 92464 0 92520 800 6 la_oen[90]
port 488 nsew signal input
rlabel metal2 s 93200 0 93256 800 6 la_oen[91]
port 489 nsew signal input
rlabel metal2 s 93936 0 93992 800 6 la_oen[92]
port 490 nsew signal input
rlabel metal2 s 94672 0 94728 800 6 la_oen[93]
port 491 nsew signal input
rlabel metal2 s 95408 0 95464 800 6 la_oen[94]
port 492 nsew signal input
rlabel metal2 s 96144 0 96200 800 6 la_oen[95]
port 493 nsew signal input
rlabel metal2 s 96880 0 96936 800 6 la_oen[96]
port 494 nsew signal input
rlabel metal2 s 97616 0 97672 800 6 la_oen[97]
port 495 nsew signal input
rlabel metal2 s 98352 0 98408 800 6 la_oen[98]
port 496 nsew signal input
rlabel metal2 s 99088 0 99144 800 6 la_oen[99]
port 497 nsew signal input
rlabel metal2 s 33032 0 33088 800 6 la_oen[9]
port 498 nsew signal input
rlabel metal2 s 4 0 60 800 6 wb_clk_i
port 499 nsew signal input
rlabel metal2 s 188 0 244 800 6 wb_rst_i
port 500 nsew signal input
rlabel metal2 s 464 0 520 800 6 wbs_ack_o
port 501 nsew signal output
rlabel metal2 s 1384 0 1440 800 6 wbs_adr_i[0]
port 502 nsew signal input
rlabel metal2 s 9756 0 9812 800 6 wbs_adr_i[10]
port 503 nsew signal input
rlabel metal2 s 10492 0 10548 800 6 wbs_adr_i[11]
port 504 nsew signal input
rlabel metal2 s 11228 0 11284 800 6 wbs_adr_i[12]
port 505 nsew signal input
rlabel metal2 s 11964 0 12020 800 6 wbs_adr_i[13]
port 506 nsew signal input
rlabel metal2 s 12700 0 12756 800 6 wbs_adr_i[14]
port 507 nsew signal input
rlabel metal2 s 13436 0 13492 800 6 wbs_adr_i[15]
port 508 nsew signal input
rlabel metal2 s 14172 0 14228 800 6 wbs_adr_i[16]
port 509 nsew signal input
rlabel metal2 s 14908 0 14964 800 6 wbs_adr_i[17]
port 510 nsew signal input
rlabel metal2 s 15644 0 15700 800 6 wbs_adr_i[18]
port 511 nsew signal input
rlabel metal2 s 16380 0 16436 800 6 wbs_adr_i[19]
port 512 nsew signal input
rlabel metal2 s 2396 0 2452 800 6 wbs_adr_i[1]
port 513 nsew signal input
rlabel metal2 s 17116 0 17172 800 6 wbs_adr_i[20]
port 514 nsew signal input
rlabel metal2 s 17852 0 17908 800 6 wbs_adr_i[21]
port 515 nsew signal input
rlabel metal2 s 18588 0 18644 800 6 wbs_adr_i[22]
port 516 nsew signal input
rlabel metal2 s 19324 0 19380 800 6 wbs_adr_i[23]
port 517 nsew signal input
rlabel metal2 s 20060 0 20116 800 6 wbs_adr_i[24]
port 518 nsew signal input
rlabel metal2 s 20796 0 20852 800 6 wbs_adr_i[25]
port 519 nsew signal input
rlabel metal2 s 21532 0 21588 800 6 wbs_adr_i[26]
port 520 nsew signal input
rlabel metal2 s 22268 0 22324 800 6 wbs_adr_i[27]
port 521 nsew signal input
rlabel metal2 s 23004 0 23060 800 6 wbs_adr_i[28]
port 522 nsew signal input
rlabel metal2 s 23740 0 23796 800 6 wbs_adr_i[29]
port 523 nsew signal input
rlabel metal2 s 3408 0 3464 800 6 wbs_adr_i[2]
port 524 nsew signal input
rlabel metal2 s 24476 0 24532 800 6 wbs_adr_i[30]
port 525 nsew signal input
rlabel metal2 s 25212 0 25268 800 6 wbs_adr_i[31]
port 526 nsew signal input
rlabel metal2 s 4328 0 4384 800 6 wbs_adr_i[3]
port 527 nsew signal input
rlabel metal2 s 5340 0 5396 800 6 wbs_adr_i[4]
port 528 nsew signal input
rlabel metal2 s 6076 0 6132 800 6 wbs_adr_i[5]
port 529 nsew signal input
rlabel metal2 s 6812 0 6868 800 6 wbs_adr_i[6]
port 530 nsew signal input
rlabel metal2 s 7548 0 7604 800 6 wbs_adr_i[7]
port 531 nsew signal input
rlabel metal2 s 8284 0 8340 800 6 wbs_adr_i[8]
port 532 nsew signal input
rlabel metal2 s 9020 0 9076 800 6 wbs_adr_i[9]
port 533 nsew signal input
rlabel metal2 s 648 0 704 800 6 wbs_cyc_i
port 534 nsew signal input
rlabel metal2 s 1660 0 1716 800 6 wbs_dat_i[0]
port 535 nsew signal input
rlabel metal2 s 10032 0 10088 800 6 wbs_dat_i[10]
port 536 nsew signal input
rlabel metal2 s 10768 0 10824 800 6 wbs_dat_i[11]
port 537 nsew signal input
rlabel metal2 s 11504 0 11560 800 6 wbs_dat_i[12]
port 538 nsew signal input
rlabel metal2 s 12240 0 12296 800 6 wbs_dat_i[13]
port 539 nsew signal input
rlabel metal2 s 12976 0 13032 800 6 wbs_dat_i[14]
port 540 nsew signal input
rlabel metal2 s 13712 0 13768 800 6 wbs_dat_i[15]
port 541 nsew signal input
rlabel metal2 s 14448 0 14504 800 6 wbs_dat_i[16]
port 542 nsew signal input
rlabel metal2 s 15092 0 15148 800 6 wbs_dat_i[17]
port 543 nsew signal input
rlabel metal2 s 15828 0 15884 800 6 wbs_dat_i[18]
port 544 nsew signal input
rlabel metal2 s 16564 0 16620 800 6 wbs_dat_i[19]
port 545 nsew signal input
rlabel metal2 s 2672 0 2728 800 6 wbs_dat_i[1]
port 546 nsew signal input
rlabel metal2 s 17300 0 17356 800 6 wbs_dat_i[20]
port 547 nsew signal input
rlabel metal2 s 18036 0 18092 800 6 wbs_dat_i[21]
port 548 nsew signal input
rlabel metal2 s 18772 0 18828 800 6 wbs_dat_i[22]
port 549 nsew signal input
rlabel metal2 s 19508 0 19564 800 6 wbs_dat_i[23]
port 550 nsew signal input
rlabel metal2 s 20244 0 20300 800 6 wbs_dat_i[24]
port 551 nsew signal input
rlabel metal2 s 20980 0 21036 800 6 wbs_dat_i[25]
port 552 nsew signal input
rlabel metal2 s 21716 0 21772 800 6 wbs_dat_i[26]
port 553 nsew signal input
rlabel metal2 s 22452 0 22508 800 6 wbs_dat_i[27]
port 554 nsew signal input
rlabel metal2 s 23188 0 23244 800 6 wbs_dat_i[28]
port 555 nsew signal input
rlabel metal2 s 23924 0 23980 800 6 wbs_dat_i[29]
port 556 nsew signal input
rlabel metal2 s 3592 0 3648 800 6 wbs_dat_i[2]
port 557 nsew signal input
rlabel metal2 s 24660 0 24716 800 6 wbs_dat_i[30]
port 558 nsew signal input
rlabel metal2 s 25396 0 25452 800 6 wbs_dat_i[31]
port 559 nsew signal input
rlabel metal2 s 4604 0 4660 800 6 wbs_dat_i[3]
port 560 nsew signal input
rlabel metal2 s 5616 0 5672 800 6 wbs_dat_i[4]
port 561 nsew signal input
rlabel metal2 s 6352 0 6408 800 6 wbs_dat_i[5]
port 562 nsew signal input
rlabel metal2 s 7088 0 7144 800 6 wbs_dat_i[6]
port 563 nsew signal input
rlabel metal2 s 7824 0 7880 800 6 wbs_dat_i[7]
port 564 nsew signal input
rlabel metal2 s 8560 0 8616 800 6 wbs_dat_i[8]
port 565 nsew signal input
rlabel metal2 s 9296 0 9352 800 6 wbs_dat_i[9]
port 566 nsew signal input
rlabel metal2 s 1936 0 1992 800 6 wbs_dat_o[0]
port 567 nsew signal output
rlabel metal2 s 10216 0 10272 800 6 wbs_dat_o[10]
port 568 nsew signal output
rlabel metal2 s 10952 0 11008 800 6 wbs_dat_o[11]
port 569 nsew signal output
rlabel metal2 s 11688 0 11744 800 6 wbs_dat_o[12]
port 570 nsew signal output
rlabel metal2 s 12424 0 12480 800 6 wbs_dat_o[13]
port 571 nsew signal output
rlabel metal2 s 13160 0 13216 800 6 wbs_dat_o[14]
port 572 nsew signal output
rlabel metal2 s 13896 0 13952 800 6 wbs_dat_o[15]
port 573 nsew signal output
rlabel metal2 s 14632 0 14688 800 6 wbs_dat_o[16]
port 574 nsew signal output
rlabel metal2 s 15368 0 15424 800 6 wbs_dat_o[17]
port 575 nsew signal output
rlabel metal2 s 16104 0 16160 800 6 wbs_dat_o[18]
port 576 nsew signal output
rlabel metal2 s 16840 0 16896 800 6 wbs_dat_o[19]
port 577 nsew signal output
rlabel metal2 s 2856 0 2912 800 6 wbs_dat_o[1]
port 578 nsew signal output
rlabel metal2 s 17576 0 17632 800 6 wbs_dat_o[20]
port 579 nsew signal output
rlabel metal2 s 18312 0 18368 800 6 wbs_dat_o[21]
port 580 nsew signal output
rlabel metal2 s 19048 0 19104 800 6 wbs_dat_o[22]
port 581 nsew signal output
rlabel metal2 s 19784 0 19840 800 6 wbs_dat_o[23]
port 582 nsew signal output
rlabel metal2 s 20520 0 20576 800 6 wbs_dat_o[24]
port 583 nsew signal output
rlabel metal2 s 21256 0 21312 800 6 wbs_dat_o[25]
port 584 nsew signal output
rlabel metal2 s 21992 0 22048 800 6 wbs_dat_o[26]
port 585 nsew signal output
rlabel metal2 s 22728 0 22784 800 6 wbs_dat_o[27]
port 586 nsew signal output
rlabel metal2 s 23464 0 23520 800 6 wbs_dat_o[28]
port 587 nsew signal output
rlabel metal2 s 24200 0 24256 800 6 wbs_dat_o[29]
port 588 nsew signal output
rlabel metal2 s 3868 0 3924 800 6 wbs_dat_o[2]
port 589 nsew signal output
rlabel metal2 s 24936 0 24992 800 6 wbs_dat_o[30]
port 590 nsew signal output
rlabel metal2 s 25672 0 25728 800 6 wbs_dat_o[31]
port 591 nsew signal output
rlabel metal2 s 4880 0 4936 800 6 wbs_dat_o[3]
port 592 nsew signal output
rlabel metal2 s 5800 0 5856 800 6 wbs_dat_o[4]
port 593 nsew signal output
rlabel metal2 s 6536 0 6592 800 6 wbs_dat_o[5]
port 594 nsew signal output
rlabel metal2 s 7272 0 7328 800 6 wbs_dat_o[6]
port 595 nsew signal output
rlabel metal2 s 8008 0 8064 800 6 wbs_dat_o[7]
port 596 nsew signal output
rlabel metal2 s 8744 0 8800 800 6 wbs_dat_o[8]
port 597 nsew signal output
rlabel metal2 s 9480 0 9536 800 6 wbs_dat_o[9]
port 598 nsew signal output
rlabel metal2 s 2120 0 2176 800 6 wbs_sel_i[0]
port 599 nsew signal input
rlabel metal2 s 3132 0 3188 800 6 wbs_sel_i[1]
port 600 nsew signal input
rlabel metal2 s 4144 0 4200 800 6 wbs_sel_i[2]
port 601 nsew signal input
rlabel metal2 s 5064 0 5120 800 6 wbs_sel_i[3]
port 602 nsew signal input
rlabel metal2 s 924 0 980 800 6 wbs_stb_i
port 603 nsew signal input
rlabel metal2 s 1200 0 1256 800 6 wbs_we_i
port 604 nsew signal input
rlabel metal4 s 96262 2128 96582 117552 6 vccd1
port 605 nsew power bidirectional
rlabel metal4 s 65542 2128 65862 117552 6 vccd1
port 606 nsew power bidirectional
rlabel metal4 s 34822 2128 35142 117552 6 vccd1
port 607 nsew power bidirectional
rlabel metal4 s 4102 2128 4422 117552 6 vccd1
port 608 nsew power bidirectional
rlabel metal4 s 111622 2128 111942 117552 6 vssd1
port 609 nsew ground bidirectional
rlabel metal4 s 80902 2128 81222 117552 6 vssd1
port 610 nsew ground bidirectional
rlabel metal4 s 50182 2128 50502 117552 6 vssd1
port 611 nsew ground bidirectional
rlabel metal4 s 19462 2128 19782 117552 6 vssd1
port 612 nsew ground bidirectional
rlabel metal4 s 96922 2176 97242 117504 6 vccd2
port 613 nsew power bidirectional
rlabel metal4 s 66202 2176 66522 117504 6 vccd2
port 614 nsew power bidirectional
rlabel metal4 s 35482 2176 35802 117504 6 vccd2
port 615 nsew power bidirectional
rlabel metal4 s 4762 2176 5082 117504 6 vccd2
port 616 nsew power bidirectional
rlabel metal4 s 112282 2176 112602 117504 6 vssd2
port 617 nsew ground bidirectional
rlabel metal4 s 81562 2176 81882 117504 6 vssd2
port 618 nsew ground bidirectional
rlabel metal4 s 50842 2176 51162 117504 6 vssd2
port 619 nsew ground bidirectional
rlabel metal4 s 20122 2176 20442 117504 6 vssd2
port 620 nsew ground bidirectional
rlabel metal4 s 97582 2176 97902 117504 6 vdda1
port 621 nsew power bidirectional
rlabel metal4 s 66862 2176 67182 117504 6 vdda1
port 622 nsew power bidirectional
rlabel metal4 s 36142 2176 36462 117504 6 vdda1
port 623 nsew power bidirectional
rlabel metal4 s 5422 2176 5742 117504 6 vdda1
port 624 nsew power bidirectional
rlabel metal4 s 112942 2176 113262 117504 6 vssa1
port 625 nsew ground bidirectional
rlabel metal4 s 82222 2176 82542 117504 6 vssa1
port 626 nsew ground bidirectional
rlabel metal4 s 51502 2176 51822 117504 6 vssa1
port 627 nsew ground bidirectional
rlabel metal4 s 20782 2176 21102 117504 6 vssa1
port 628 nsew ground bidirectional
rlabel metal4 s 98242 2176 98562 117504 6 vdda2
port 629 nsew power bidirectional
rlabel metal4 s 67522 2176 67842 117504 6 vdda2
port 630 nsew power bidirectional
rlabel metal4 s 36802 2176 37122 117504 6 vdda2
port 631 nsew power bidirectional
rlabel metal4 s 6082 2176 6402 117504 6 vdda2
port 632 nsew power bidirectional
rlabel metal4 s 113602 2176 113922 117504 6 vssa2
port 633 nsew ground bidirectional
rlabel metal4 s 82882 2176 83202 117504 6 vssa2
port 634 nsew ground bidirectional
rlabel metal4 s 52162 2176 52482 117504 6 vssa2
port 635 nsew ground bidirectional
rlabel metal4 s 21442 2176 21762 117504 6 vssa2
port 636 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 119752 120000
string LEFview TRUE
<< end >>
